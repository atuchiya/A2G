magic
tech sky130A
magscale 1 2
timestamp 1686266350
<< checkpaint >>
rect -1899 -1619 1899 1619
<< pwell >>
rect -639 -359 639 359
<< nmos >>
rect -443 -211 -383 149
rect -325 -211 -265 149
rect -207 -211 -147 149
rect -89 -211 -29 149
rect 29 -211 89 149
rect 147 -211 207 149
rect 265 -211 325 149
rect 383 -211 443 149
<< ndiff >>
rect -501 137 -443 149
rect -501 -199 -489 137
rect -455 -199 -443 137
rect -501 -211 -443 -199
rect -383 137 -325 149
rect -383 -199 -371 137
rect -337 -199 -325 137
rect -383 -211 -325 -199
rect -265 137 -207 149
rect -265 -199 -253 137
rect -219 -199 -207 137
rect -265 -211 -207 -199
rect -147 137 -89 149
rect -147 -199 -135 137
rect -101 -199 -89 137
rect -147 -211 -89 -199
rect -29 137 29 149
rect -29 -199 -17 137
rect 17 -199 29 137
rect -29 -211 29 -199
rect 89 137 147 149
rect 89 -199 101 137
rect 135 -199 147 137
rect 89 -211 147 -199
rect 207 137 265 149
rect 207 -199 219 137
rect 253 -199 265 137
rect 207 -211 265 -199
rect 325 137 383 149
rect 325 -199 337 137
rect 371 -199 383 137
rect 325 -211 383 -199
rect 443 137 501 149
rect 443 -199 455 137
rect 489 -199 501 137
rect 443 -211 501 -199
<< ndiffc >>
rect -489 -199 -455 137
rect -371 -199 -337 137
rect -253 -199 -219 137
rect -135 -199 -101 137
rect -17 -199 17 137
rect 101 -199 135 137
rect 219 -199 253 137
rect 337 -199 371 137
rect 455 -199 489 137
<< psubdiff >>
rect -603 289 -507 323
rect 507 289 603 323
rect -603 227 -569 289
rect 569 227 603 289
rect -603 -289 -569 -227
rect 569 -289 603 -227
rect -603 -323 -507 -289
rect 507 -323 603 -289
<< psubdiffcont >>
rect -507 289 507 323
rect -603 -227 -569 227
rect 569 -227 603 227
rect -507 -323 507 -289
<< poly >>
rect -446 221 -380 237
rect -446 187 -430 221
rect -396 187 -380 221
rect -446 171 -380 187
rect -328 221 -262 237
rect -328 187 -312 221
rect -278 187 -262 221
rect -328 171 -262 187
rect -210 221 -144 237
rect -210 187 -194 221
rect -160 187 -144 221
rect -210 171 -144 187
rect -92 221 -26 237
rect -92 187 -76 221
rect -42 187 -26 221
rect -92 171 -26 187
rect 26 221 92 237
rect 26 187 42 221
rect 76 187 92 221
rect 26 171 92 187
rect 144 221 210 237
rect 144 187 160 221
rect 194 187 210 221
rect 144 171 210 187
rect 262 221 328 237
rect 262 187 278 221
rect 312 187 328 221
rect 262 171 328 187
rect 380 221 446 237
rect 380 187 396 221
rect 430 187 446 221
rect 380 171 446 187
rect -443 149 -383 171
rect -325 149 -265 171
rect -207 149 -147 171
rect -89 149 -29 171
rect 29 149 89 171
rect 147 149 207 171
rect 265 149 325 171
rect 383 149 443 171
rect -443 -237 -383 -211
rect -325 -237 -265 -211
rect -207 -237 -147 -211
rect -89 -237 -29 -211
rect 29 -237 89 -211
rect 147 -237 207 -211
rect 265 -237 325 -211
rect 383 -237 443 -211
<< polycont >>
rect -430 187 -396 221
rect -312 187 -278 221
rect -194 187 -160 221
rect -76 187 -42 221
rect 42 187 76 221
rect 160 187 194 221
rect 278 187 312 221
rect 396 187 430 221
<< locali >>
rect -603 289 -507 323
rect 507 289 603 323
rect -603 227 -569 289
rect 569 227 603 289
rect -446 187 -430 221
rect -396 187 -380 221
rect -328 187 -312 221
rect -278 187 -262 221
rect -210 187 -194 221
rect -160 187 -144 221
rect -92 187 -76 221
rect -42 187 -26 221
rect 26 187 42 221
rect 76 187 92 221
rect 144 187 160 221
rect 194 187 210 221
rect 262 187 278 221
rect 312 187 328 221
rect 380 187 396 221
rect 430 187 446 221
rect -489 137 -455 153
rect -489 -215 -455 -199
rect -371 137 -337 153
rect -371 -215 -337 -199
rect -253 137 -219 153
rect -253 -215 -219 -199
rect -135 137 -101 153
rect -135 -215 -101 -199
rect -17 137 17 153
rect -17 -215 17 -199
rect 101 137 135 153
rect 101 -215 135 -199
rect 219 137 253 153
rect 219 -215 253 -199
rect 337 137 371 153
rect 337 -215 371 -199
rect 455 137 489 153
rect 455 -215 489 -199
rect -603 -289 -569 -227
rect 569 -289 603 -227
rect -603 -323 -507 -289
rect 507 -323 603 -289
<< viali >>
rect -430 187 -396 221
rect -312 187 -278 221
rect -194 187 -160 221
rect -76 187 -42 221
rect 42 187 76 221
rect 160 187 194 221
rect 278 187 312 221
rect 396 187 430 221
rect -489 -199 -455 137
rect -371 -199 -337 137
rect -253 -199 -219 137
rect -135 -199 -101 137
rect -17 -199 17 137
rect 101 -199 135 137
rect 219 -199 253 137
rect 337 -199 371 137
rect 455 -199 489 137
<< metal1 >>
rect -442 221 -384 227
rect -442 187 -430 221
rect -396 187 -384 221
rect -442 181 -384 187
rect -324 221 -266 227
rect -324 187 -312 221
rect -278 187 -266 221
rect -324 181 -266 187
rect -206 221 -148 227
rect -206 187 -194 221
rect -160 187 -148 221
rect -206 181 -148 187
rect -88 221 -30 227
rect -88 187 -76 221
rect -42 187 -30 221
rect -88 181 -30 187
rect 30 221 88 227
rect 30 187 42 221
rect 76 187 88 221
rect 30 181 88 187
rect 148 221 206 227
rect 148 187 160 221
rect 194 187 206 221
rect 148 181 206 187
rect 266 221 324 227
rect 266 187 278 221
rect 312 187 324 221
rect 266 181 324 187
rect 384 221 442 227
rect 384 187 396 221
rect 430 187 442 221
rect 384 181 442 187
rect -495 137 -449 149
rect -495 -199 -489 137
rect -455 -199 -449 137
rect -495 -211 -449 -199
rect -377 137 -331 149
rect -377 -199 -371 137
rect -337 -199 -331 137
rect -377 -211 -331 -199
rect -259 137 -213 149
rect -259 -199 -253 137
rect -219 -199 -213 137
rect -259 -211 -213 -199
rect -141 137 -95 149
rect -141 -199 -135 137
rect -101 -199 -95 137
rect -141 -211 -95 -199
rect -23 137 23 149
rect -23 -199 -17 137
rect 17 -199 23 137
rect -23 -211 23 -199
rect 95 137 141 149
rect 95 -199 101 137
rect 135 -199 141 137
rect 95 -211 141 -199
rect 213 137 259 149
rect 213 -199 219 137
rect 253 -199 259 137
rect 213 -211 259 -199
rect 331 137 377 149
rect 331 -199 337 137
rect 371 -199 377 137
rect 331 -211 377 -199
rect 449 137 495 149
rect 449 -199 455 137
rect 489 -199 495 137
rect 449 -211 495 -199
<< labels >>
flabel metal1 -413 204 -413 204 0 FreeSans 240 0 0 0 G
flabel metal1 -295 204 -295 204 0 FreeSans 240 0 0 0 G
flabel metal1 -177 204 -177 204 0 FreeSans 240 0 0 0 G
flabel metal1 -59 204 -59 204 0 FreeSans 240 0 0 0 G
flabel metal1 59 204 59 204 0 FreeSans 240 0 0 0 G
flabel metal1 177 204 177 204 0 FreeSans 240 0 0 0 G
flabel metal1 295 204 295 204 0 FreeSans 240 0 0 0 G
flabel metal1 413 204 413 204 0 FreeSans 240 0 0 0 G
flabel metal1 -472 -31 -472 -31 0 FreeSans 240 0 0 0 D
flabel metal1 -354 -31 -354 -31 0 FreeSans 240 0 0 0 S
flabel metal1 -236 -31 -236 -31 0 FreeSans 240 0 0 0 D
flabel metal1 -118 -31 -118 -31 0 FreeSans 240 0 0 0 S
flabel metal1 0 -31 0 -31 0 FreeSans 240 0 0 0 D
flabel metal1 118 -31 118 -31 0 FreeSans 240 0 0 0 S
flabel metal1 236 -31 236 -31 0 FreeSans 240 0 0 0 D
flabel metal1 354 -31 354 -31 0 FreeSans 240 0 0 0 S
flabel metal1 472 -31 472 -31 0 FreeSans 240 0 0 0 D
<< properties >>
string FIXED_BBOX -586 -306 586 306
<< end >>

