magic
tech sky130A
magscale 1 2
timestamp 1680002671
<< error_p >>
rect -2527 395 -2465 401
rect -2399 395 -2337 401
rect -2271 395 -2209 401
rect -2143 395 -2081 401
rect -2015 395 -1953 401
rect -1887 395 -1825 401
rect -1759 395 -1697 401
rect -1631 395 -1569 401
rect -1503 395 -1441 401
rect -1375 395 -1313 401
rect -1247 395 -1185 401
rect -1119 395 -1057 401
rect -991 395 -929 401
rect -863 395 -801 401
rect -735 395 -673 401
rect -607 395 -545 401
rect -479 395 -417 401
rect -351 395 -289 401
rect -223 395 -161 401
rect -95 395 -33 401
rect 33 395 95 401
rect 161 395 223 401
rect 289 395 351 401
rect 417 395 479 401
rect 545 395 607 401
rect 673 395 735 401
rect 801 395 863 401
rect 929 395 991 401
rect 1057 395 1119 401
rect 1185 395 1247 401
rect 1313 395 1375 401
rect 1441 395 1503 401
rect 1569 395 1631 401
rect 1697 395 1759 401
rect 1825 395 1887 401
rect 1953 395 2015 401
rect 2081 395 2143 401
rect 2209 395 2271 401
rect 2337 395 2399 401
rect 2465 395 2527 401
rect -2527 361 -2513 395
rect -2399 361 -2385 395
rect -2271 361 -2257 395
rect -2143 361 -2129 395
rect -2015 361 -2001 395
rect -1887 361 -1873 395
rect -1759 361 -1745 395
rect -1631 361 -1617 395
rect -1503 361 -1489 395
rect -1375 361 -1361 395
rect -1247 361 -1233 395
rect -1119 361 -1105 395
rect -991 361 -977 395
rect -863 361 -849 395
rect -735 361 -721 395
rect -607 361 -593 395
rect -479 361 -465 395
rect -351 361 -337 395
rect -223 361 -209 395
rect -95 361 -81 395
rect 33 361 47 395
rect 161 361 175 395
rect 289 361 303 395
rect 417 361 431 395
rect 545 361 559 395
rect 673 361 687 395
rect 801 361 815 395
rect 929 361 943 395
rect 1057 361 1071 395
rect 1185 361 1199 395
rect 1313 361 1327 395
rect 1441 361 1455 395
rect 1569 361 1583 395
rect 1697 361 1711 395
rect 1825 361 1839 395
rect 1953 361 1967 395
rect 2081 361 2095 395
rect 2209 361 2223 395
rect 2337 361 2351 395
rect 2465 361 2479 395
rect -2527 355 -2465 361
rect -2399 355 -2337 361
rect -2271 355 -2209 361
rect -2143 355 -2081 361
rect -2015 355 -1953 361
rect -1887 355 -1825 361
rect -1759 355 -1697 361
rect -1631 355 -1569 361
rect -1503 355 -1441 361
rect -1375 355 -1313 361
rect -1247 355 -1185 361
rect -1119 355 -1057 361
rect -991 355 -929 361
rect -863 355 -801 361
rect -735 355 -673 361
rect -607 355 -545 361
rect -479 355 -417 361
rect -351 355 -289 361
rect -223 355 -161 361
rect -95 355 -33 361
rect 33 355 95 361
rect 161 355 223 361
rect 289 355 351 361
rect 417 355 479 361
rect 545 355 607 361
rect 673 355 735 361
rect 801 355 863 361
rect 929 355 991 361
rect 1057 355 1119 361
rect 1185 355 1247 361
rect 1313 355 1375 361
rect 1441 355 1503 361
rect 1569 355 1631 361
rect 1697 355 1759 361
rect 1825 355 1887 361
rect 1953 355 2015 361
rect 2081 355 2143 361
rect 2209 355 2271 361
rect 2337 355 2399 361
rect 2465 355 2527 361
<< nwell >>
rect -2727 -534 2727 534
<< pmoslvt >>
rect -2531 -386 -2461 314
rect -2403 -386 -2333 314
rect -2275 -386 -2205 314
rect -2147 -386 -2077 314
rect -2019 -386 -1949 314
rect -1891 -386 -1821 314
rect -1763 -386 -1693 314
rect -1635 -386 -1565 314
rect -1507 -386 -1437 314
rect -1379 -386 -1309 314
rect -1251 -386 -1181 314
rect -1123 -386 -1053 314
rect -995 -386 -925 314
rect -867 -386 -797 314
rect -739 -386 -669 314
rect -611 -386 -541 314
rect -483 -386 -413 314
rect -355 -386 -285 314
rect -227 -386 -157 314
rect -99 -386 -29 314
rect 29 -386 99 314
rect 157 -386 227 314
rect 285 -386 355 314
rect 413 -386 483 314
rect 541 -386 611 314
rect 669 -386 739 314
rect 797 -386 867 314
rect 925 -386 995 314
rect 1053 -386 1123 314
rect 1181 -386 1251 314
rect 1309 -386 1379 314
rect 1437 -386 1507 314
rect 1565 -386 1635 314
rect 1693 -386 1763 314
rect 1821 -386 1891 314
rect 1949 -386 2019 314
rect 2077 -386 2147 314
rect 2205 -386 2275 314
rect 2333 -386 2403 314
rect 2461 -386 2531 314
<< pdiff >>
rect -2589 287 -2531 314
rect -2589 253 -2577 287
rect -2543 253 -2531 287
rect -2589 219 -2531 253
rect -2589 185 -2577 219
rect -2543 185 -2531 219
rect -2589 151 -2531 185
rect -2589 117 -2577 151
rect -2543 117 -2531 151
rect -2589 83 -2531 117
rect -2589 49 -2577 83
rect -2543 49 -2531 83
rect -2589 15 -2531 49
rect -2589 -19 -2577 15
rect -2543 -19 -2531 15
rect -2589 -53 -2531 -19
rect -2589 -87 -2577 -53
rect -2543 -87 -2531 -53
rect -2589 -121 -2531 -87
rect -2589 -155 -2577 -121
rect -2543 -155 -2531 -121
rect -2589 -189 -2531 -155
rect -2589 -223 -2577 -189
rect -2543 -223 -2531 -189
rect -2589 -257 -2531 -223
rect -2589 -291 -2577 -257
rect -2543 -291 -2531 -257
rect -2589 -325 -2531 -291
rect -2589 -359 -2577 -325
rect -2543 -359 -2531 -325
rect -2589 -386 -2531 -359
rect -2461 287 -2403 314
rect -2461 253 -2449 287
rect -2415 253 -2403 287
rect -2461 219 -2403 253
rect -2461 185 -2449 219
rect -2415 185 -2403 219
rect -2461 151 -2403 185
rect -2461 117 -2449 151
rect -2415 117 -2403 151
rect -2461 83 -2403 117
rect -2461 49 -2449 83
rect -2415 49 -2403 83
rect -2461 15 -2403 49
rect -2461 -19 -2449 15
rect -2415 -19 -2403 15
rect -2461 -53 -2403 -19
rect -2461 -87 -2449 -53
rect -2415 -87 -2403 -53
rect -2461 -121 -2403 -87
rect -2461 -155 -2449 -121
rect -2415 -155 -2403 -121
rect -2461 -189 -2403 -155
rect -2461 -223 -2449 -189
rect -2415 -223 -2403 -189
rect -2461 -257 -2403 -223
rect -2461 -291 -2449 -257
rect -2415 -291 -2403 -257
rect -2461 -325 -2403 -291
rect -2461 -359 -2449 -325
rect -2415 -359 -2403 -325
rect -2461 -386 -2403 -359
rect -2333 287 -2275 314
rect -2333 253 -2321 287
rect -2287 253 -2275 287
rect -2333 219 -2275 253
rect -2333 185 -2321 219
rect -2287 185 -2275 219
rect -2333 151 -2275 185
rect -2333 117 -2321 151
rect -2287 117 -2275 151
rect -2333 83 -2275 117
rect -2333 49 -2321 83
rect -2287 49 -2275 83
rect -2333 15 -2275 49
rect -2333 -19 -2321 15
rect -2287 -19 -2275 15
rect -2333 -53 -2275 -19
rect -2333 -87 -2321 -53
rect -2287 -87 -2275 -53
rect -2333 -121 -2275 -87
rect -2333 -155 -2321 -121
rect -2287 -155 -2275 -121
rect -2333 -189 -2275 -155
rect -2333 -223 -2321 -189
rect -2287 -223 -2275 -189
rect -2333 -257 -2275 -223
rect -2333 -291 -2321 -257
rect -2287 -291 -2275 -257
rect -2333 -325 -2275 -291
rect -2333 -359 -2321 -325
rect -2287 -359 -2275 -325
rect -2333 -386 -2275 -359
rect -2205 287 -2147 314
rect -2205 253 -2193 287
rect -2159 253 -2147 287
rect -2205 219 -2147 253
rect -2205 185 -2193 219
rect -2159 185 -2147 219
rect -2205 151 -2147 185
rect -2205 117 -2193 151
rect -2159 117 -2147 151
rect -2205 83 -2147 117
rect -2205 49 -2193 83
rect -2159 49 -2147 83
rect -2205 15 -2147 49
rect -2205 -19 -2193 15
rect -2159 -19 -2147 15
rect -2205 -53 -2147 -19
rect -2205 -87 -2193 -53
rect -2159 -87 -2147 -53
rect -2205 -121 -2147 -87
rect -2205 -155 -2193 -121
rect -2159 -155 -2147 -121
rect -2205 -189 -2147 -155
rect -2205 -223 -2193 -189
rect -2159 -223 -2147 -189
rect -2205 -257 -2147 -223
rect -2205 -291 -2193 -257
rect -2159 -291 -2147 -257
rect -2205 -325 -2147 -291
rect -2205 -359 -2193 -325
rect -2159 -359 -2147 -325
rect -2205 -386 -2147 -359
rect -2077 287 -2019 314
rect -2077 253 -2065 287
rect -2031 253 -2019 287
rect -2077 219 -2019 253
rect -2077 185 -2065 219
rect -2031 185 -2019 219
rect -2077 151 -2019 185
rect -2077 117 -2065 151
rect -2031 117 -2019 151
rect -2077 83 -2019 117
rect -2077 49 -2065 83
rect -2031 49 -2019 83
rect -2077 15 -2019 49
rect -2077 -19 -2065 15
rect -2031 -19 -2019 15
rect -2077 -53 -2019 -19
rect -2077 -87 -2065 -53
rect -2031 -87 -2019 -53
rect -2077 -121 -2019 -87
rect -2077 -155 -2065 -121
rect -2031 -155 -2019 -121
rect -2077 -189 -2019 -155
rect -2077 -223 -2065 -189
rect -2031 -223 -2019 -189
rect -2077 -257 -2019 -223
rect -2077 -291 -2065 -257
rect -2031 -291 -2019 -257
rect -2077 -325 -2019 -291
rect -2077 -359 -2065 -325
rect -2031 -359 -2019 -325
rect -2077 -386 -2019 -359
rect -1949 287 -1891 314
rect -1949 253 -1937 287
rect -1903 253 -1891 287
rect -1949 219 -1891 253
rect -1949 185 -1937 219
rect -1903 185 -1891 219
rect -1949 151 -1891 185
rect -1949 117 -1937 151
rect -1903 117 -1891 151
rect -1949 83 -1891 117
rect -1949 49 -1937 83
rect -1903 49 -1891 83
rect -1949 15 -1891 49
rect -1949 -19 -1937 15
rect -1903 -19 -1891 15
rect -1949 -53 -1891 -19
rect -1949 -87 -1937 -53
rect -1903 -87 -1891 -53
rect -1949 -121 -1891 -87
rect -1949 -155 -1937 -121
rect -1903 -155 -1891 -121
rect -1949 -189 -1891 -155
rect -1949 -223 -1937 -189
rect -1903 -223 -1891 -189
rect -1949 -257 -1891 -223
rect -1949 -291 -1937 -257
rect -1903 -291 -1891 -257
rect -1949 -325 -1891 -291
rect -1949 -359 -1937 -325
rect -1903 -359 -1891 -325
rect -1949 -386 -1891 -359
rect -1821 287 -1763 314
rect -1821 253 -1809 287
rect -1775 253 -1763 287
rect -1821 219 -1763 253
rect -1821 185 -1809 219
rect -1775 185 -1763 219
rect -1821 151 -1763 185
rect -1821 117 -1809 151
rect -1775 117 -1763 151
rect -1821 83 -1763 117
rect -1821 49 -1809 83
rect -1775 49 -1763 83
rect -1821 15 -1763 49
rect -1821 -19 -1809 15
rect -1775 -19 -1763 15
rect -1821 -53 -1763 -19
rect -1821 -87 -1809 -53
rect -1775 -87 -1763 -53
rect -1821 -121 -1763 -87
rect -1821 -155 -1809 -121
rect -1775 -155 -1763 -121
rect -1821 -189 -1763 -155
rect -1821 -223 -1809 -189
rect -1775 -223 -1763 -189
rect -1821 -257 -1763 -223
rect -1821 -291 -1809 -257
rect -1775 -291 -1763 -257
rect -1821 -325 -1763 -291
rect -1821 -359 -1809 -325
rect -1775 -359 -1763 -325
rect -1821 -386 -1763 -359
rect -1693 287 -1635 314
rect -1693 253 -1681 287
rect -1647 253 -1635 287
rect -1693 219 -1635 253
rect -1693 185 -1681 219
rect -1647 185 -1635 219
rect -1693 151 -1635 185
rect -1693 117 -1681 151
rect -1647 117 -1635 151
rect -1693 83 -1635 117
rect -1693 49 -1681 83
rect -1647 49 -1635 83
rect -1693 15 -1635 49
rect -1693 -19 -1681 15
rect -1647 -19 -1635 15
rect -1693 -53 -1635 -19
rect -1693 -87 -1681 -53
rect -1647 -87 -1635 -53
rect -1693 -121 -1635 -87
rect -1693 -155 -1681 -121
rect -1647 -155 -1635 -121
rect -1693 -189 -1635 -155
rect -1693 -223 -1681 -189
rect -1647 -223 -1635 -189
rect -1693 -257 -1635 -223
rect -1693 -291 -1681 -257
rect -1647 -291 -1635 -257
rect -1693 -325 -1635 -291
rect -1693 -359 -1681 -325
rect -1647 -359 -1635 -325
rect -1693 -386 -1635 -359
rect -1565 287 -1507 314
rect -1565 253 -1553 287
rect -1519 253 -1507 287
rect -1565 219 -1507 253
rect -1565 185 -1553 219
rect -1519 185 -1507 219
rect -1565 151 -1507 185
rect -1565 117 -1553 151
rect -1519 117 -1507 151
rect -1565 83 -1507 117
rect -1565 49 -1553 83
rect -1519 49 -1507 83
rect -1565 15 -1507 49
rect -1565 -19 -1553 15
rect -1519 -19 -1507 15
rect -1565 -53 -1507 -19
rect -1565 -87 -1553 -53
rect -1519 -87 -1507 -53
rect -1565 -121 -1507 -87
rect -1565 -155 -1553 -121
rect -1519 -155 -1507 -121
rect -1565 -189 -1507 -155
rect -1565 -223 -1553 -189
rect -1519 -223 -1507 -189
rect -1565 -257 -1507 -223
rect -1565 -291 -1553 -257
rect -1519 -291 -1507 -257
rect -1565 -325 -1507 -291
rect -1565 -359 -1553 -325
rect -1519 -359 -1507 -325
rect -1565 -386 -1507 -359
rect -1437 287 -1379 314
rect -1437 253 -1425 287
rect -1391 253 -1379 287
rect -1437 219 -1379 253
rect -1437 185 -1425 219
rect -1391 185 -1379 219
rect -1437 151 -1379 185
rect -1437 117 -1425 151
rect -1391 117 -1379 151
rect -1437 83 -1379 117
rect -1437 49 -1425 83
rect -1391 49 -1379 83
rect -1437 15 -1379 49
rect -1437 -19 -1425 15
rect -1391 -19 -1379 15
rect -1437 -53 -1379 -19
rect -1437 -87 -1425 -53
rect -1391 -87 -1379 -53
rect -1437 -121 -1379 -87
rect -1437 -155 -1425 -121
rect -1391 -155 -1379 -121
rect -1437 -189 -1379 -155
rect -1437 -223 -1425 -189
rect -1391 -223 -1379 -189
rect -1437 -257 -1379 -223
rect -1437 -291 -1425 -257
rect -1391 -291 -1379 -257
rect -1437 -325 -1379 -291
rect -1437 -359 -1425 -325
rect -1391 -359 -1379 -325
rect -1437 -386 -1379 -359
rect -1309 287 -1251 314
rect -1309 253 -1297 287
rect -1263 253 -1251 287
rect -1309 219 -1251 253
rect -1309 185 -1297 219
rect -1263 185 -1251 219
rect -1309 151 -1251 185
rect -1309 117 -1297 151
rect -1263 117 -1251 151
rect -1309 83 -1251 117
rect -1309 49 -1297 83
rect -1263 49 -1251 83
rect -1309 15 -1251 49
rect -1309 -19 -1297 15
rect -1263 -19 -1251 15
rect -1309 -53 -1251 -19
rect -1309 -87 -1297 -53
rect -1263 -87 -1251 -53
rect -1309 -121 -1251 -87
rect -1309 -155 -1297 -121
rect -1263 -155 -1251 -121
rect -1309 -189 -1251 -155
rect -1309 -223 -1297 -189
rect -1263 -223 -1251 -189
rect -1309 -257 -1251 -223
rect -1309 -291 -1297 -257
rect -1263 -291 -1251 -257
rect -1309 -325 -1251 -291
rect -1309 -359 -1297 -325
rect -1263 -359 -1251 -325
rect -1309 -386 -1251 -359
rect -1181 287 -1123 314
rect -1181 253 -1169 287
rect -1135 253 -1123 287
rect -1181 219 -1123 253
rect -1181 185 -1169 219
rect -1135 185 -1123 219
rect -1181 151 -1123 185
rect -1181 117 -1169 151
rect -1135 117 -1123 151
rect -1181 83 -1123 117
rect -1181 49 -1169 83
rect -1135 49 -1123 83
rect -1181 15 -1123 49
rect -1181 -19 -1169 15
rect -1135 -19 -1123 15
rect -1181 -53 -1123 -19
rect -1181 -87 -1169 -53
rect -1135 -87 -1123 -53
rect -1181 -121 -1123 -87
rect -1181 -155 -1169 -121
rect -1135 -155 -1123 -121
rect -1181 -189 -1123 -155
rect -1181 -223 -1169 -189
rect -1135 -223 -1123 -189
rect -1181 -257 -1123 -223
rect -1181 -291 -1169 -257
rect -1135 -291 -1123 -257
rect -1181 -325 -1123 -291
rect -1181 -359 -1169 -325
rect -1135 -359 -1123 -325
rect -1181 -386 -1123 -359
rect -1053 287 -995 314
rect -1053 253 -1041 287
rect -1007 253 -995 287
rect -1053 219 -995 253
rect -1053 185 -1041 219
rect -1007 185 -995 219
rect -1053 151 -995 185
rect -1053 117 -1041 151
rect -1007 117 -995 151
rect -1053 83 -995 117
rect -1053 49 -1041 83
rect -1007 49 -995 83
rect -1053 15 -995 49
rect -1053 -19 -1041 15
rect -1007 -19 -995 15
rect -1053 -53 -995 -19
rect -1053 -87 -1041 -53
rect -1007 -87 -995 -53
rect -1053 -121 -995 -87
rect -1053 -155 -1041 -121
rect -1007 -155 -995 -121
rect -1053 -189 -995 -155
rect -1053 -223 -1041 -189
rect -1007 -223 -995 -189
rect -1053 -257 -995 -223
rect -1053 -291 -1041 -257
rect -1007 -291 -995 -257
rect -1053 -325 -995 -291
rect -1053 -359 -1041 -325
rect -1007 -359 -995 -325
rect -1053 -386 -995 -359
rect -925 287 -867 314
rect -925 253 -913 287
rect -879 253 -867 287
rect -925 219 -867 253
rect -925 185 -913 219
rect -879 185 -867 219
rect -925 151 -867 185
rect -925 117 -913 151
rect -879 117 -867 151
rect -925 83 -867 117
rect -925 49 -913 83
rect -879 49 -867 83
rect -925 15 -867 49
rect -925 -19 -913 15
rect -879 -19 -867 15
rect -925 -53 -867 -19
rect -925 -87 -913 -53
rect -879 -87 -867 -53
rect -925 -121 -867 -87
rect -925 -155 -913 -121
rect -879 -155 -867 -121
rect -925 -189 -867 -155
rect -925 -223 -913 -189
rect -879 -223 -867 -189
rect -925 -257 -867 -223
rect -925 -291 -913 -257
rect -879 -291 -867 -257
rect -925 -325 -867 -291
rect -925 -359 -913 -325
rect -879 -359 -867 -325
rect -925 -386 -867 -359
rect -797 287 -739 314
rect -797 253 -785 287
rect -751 253 -739 287
rect -797 219 -739 253
rect -797 185 -785 219
rect -751 185 -739 219
rect -797 151 -739 185
rect -797 117 -785 151
rect -751 117 -739 151
rect -797 83 -739 117
rect -797 49 -785 83
rect -751 49 -739 83
rect -797 15 -739 49
rect -797 -19 -785 15
rect -751 -19 -739 15
rect -797 -53 -739 -19
rect -797 -87 -785 -53
rect -751 -87 -739 -53
rect -797 -121 -739 -87
rect -797 -155 -785 -121
rect -751 -155 -739 -121
rect -797 -189 -739 -155
rect -797 -223 -785 -189
rect -751 -223 -739 -189
rect -797 -257 -739 -223
rect -797 -291 -785 -257
rect -751 -291 -739 -257
rect -797 -325 -739 -291
rect -797 -359 -785 -325
rect -751 -359 -739 -325
rect -797 -386 -739 -359
rect -669 287 -611 314
rect -669 253 -657 287
rect -623 253 -611 287
rect -669 219 -611 253
rect -669 185 -657 219
rect -623 185 -611 219
rect -669 151 -611 185
rect -669 117 -657 151
rect -623 117 -611 151
rect -669 83 -611 117
rect -669 49 -657 83
rect -623 49 -611 83
rect -669 15 -611 49
rect -669 -19 -657 15
rect -623 -19 -611 15
rect -669 -53 -611 -19
rect -669 -87 -657 -53
rect -623 -87 -611 -53
rect -669 -121 -611 -87
rect -669 -155 -657 -121
rect -623 -155 -611 -121
rect -669 -189 -611 -155
rect -669 -223 -657 -189
rect -623 -223 -611 -189
rect -669 -257 -611 -223
rect -669 -291 -657 -257
rect -623 -291 -611 -257
rect -669 -325 -611 -291
rect -669 -359 -657 -325
rect -623 -359 -611 -325
rect -669 -386 -611 -359
rect -541 287 -483 314
rect -541 253 -529 287
rect -495 253 -483 287
rect -541 219 -483 253
rect -541 185 -529 219
rect -495 185 -483 219
rect -541 151 -483 185
rect -541 117 -529 151
rect -495 117 -483 151
rect -541 83 -483 117
rect -541 49 -529 83
rect -495 49 -483 83
rect -541 15 -483 49
rect -541 -19 -529 15
rect -495 -19 -483 15
rect -541 -53 -483 -19
rect -541 -87 -529 -53
rect -495 -87 -483 -53
rect -541 -121 -483 -87
rect -541 -155 -529 -121
rect -495 -155 -483 -121
rect -541 -189 -483 -155
rect -541 -223 -529 -189
rect -495 -223 -483 -189
rect -541 -257 -483 -223
rect -541 -291 -529 -257
rect -495 -291 -483 -257
rect -541 -325 -483 -291
rect -541 -359 -529 -325
rect -495 -359 -483 -325
rect -541 -386 -483 -359
rect -413 287 -355 314
rect -413 253 -401 287
rect -367 253 -355 287
rect -413 219 -355 253
rect -413 185 -401 219
rect -367 185 -355 219
rect -413 151 -355 185
rect -413 117 -401 151
rect -367 117 -355 151
rect -413 83 -355 117
rect -413 49 -401 83
rect -367 49 -355 83
rect -413 15 -355 49
rect -413 -19 -401 15
rect -367 -19 -355 15
rect -413 -53 -355 -19
rect -413 -87 -401 -53
rect -367 -87 -355 -53
rect -413 -121 -355 -87
rect -413 -155 -401 -121
rect -367 -155 -355 -121
rect -413 -189 -355 -155
rect -413 -223 -401 -189
rect -367 -223 -355 -189
rect -413 -257 -355 -223
rect -413 -291 -401 -257
rect -367 -291 -355 -257
rect -413 -325 -355 -291
rect -413 -359 -401 -325
rect -367 -359 -355 -325
rect -413 -386 -355 -359
rect -285 287 -227 314
rect -285 253 -273 287
rect -239 253 -227 287
rect -285 219 -227 253
rect -285 185 -273 219
rect -239 185 -227 219
rect -285 151 -227 185
rect -285 117 -273 151
rect -239 117 -227 151
rect -285 83 -227 117
rect -285 49 -273 83
rect -239 49 -227 83
rect -285 15 -227 49
rect -285 -19 -273 15
rect -239 -19 -227 15
rect -285 -53 -227 -19
rect -285 -87 -273 -53
rect -239 -87 -227 -53
rect -285 -121 -227 -87
rect -285 -155 -273 -121
rect -239 -155 -227 -121
rect -285 -189 -227 -155
rect -285 -223 -273 -189
rect -239 -223 -227 -189
rect -285 -257 -227 -223
rect -285 -291 -273 -257
rect -239 -291 -227 -257
rect -285 -325 -227 -291
rect -285 -359 -273 -325
rect -239 -359 -227 -325
rect -285 -386 -227 -359
rect -157 287 -99 314
rect -157 253 -145 287
rect -111 253 -99 287
rect -157 219 -99 253
rect -157 185 -145 219
rect -111 185 -99 219
rect -157 151 -99 185
rect -157 117 -145 151
rect -111 117 -99 151
rect -157 83 -99 117
rect -157 49 -145 83
rect -111 49 -99 83
rect -157 15 -99 49
rect -157 -19 -145 15
rect -111 -19 -99 15
rect -157 -53 -99 -19
rect -157 -87 -145 -53
rect -111 -87 -99 -53
rect -157 -121 -99 -87
rect -157 -155 -145 -121
rect -111 -155 -99 -121
rect -157 -189 -99 -155
rect -157 -223 -145 -189
rect -111 -223 -99 -189
rect -157 -257 -99 -223
rect -157 -291 -145 -257
rect -111 -291 -99 -257
rect -157 -325 -99 -291
rect -157 -359 -145 -325
rect -111 -359 -99 -325
rect -157 -386 -99 -359
rect -29 287 29 314
rect -29 253 -17 287
rect 17 253 29 287
rect -29 219 29 253
rect -29 185 -17 219
rect 17 185 29 219
rect -29 151 29 185
rect -29 117 -17 151
rect 17 117 29 151
rect -29 83 29 117
rect -29 49 -17 83
rect 17 49 29 83
rect -29 15 29 49
rect -29 -19 -17 15
rect 17 -19 29 15
rect -29 -53 29 -19
rect -29 -87 -17 -53
rect 17 -87 29 -53
rect -29 -121 29 -87
rect -29 -155 -17 -121
rect 17 -155 29 -121
rect -29 -189 29 -155
rect -29 -223 -17 -189
rect 17 -223 29 -189
rect -29 -257 29 -223
rect -29 -291 -17 -257
rect 17 -291 29 -257
rect -29 -325 29 -291
rect -29 -359 -17 -325
rect 17 -359 29 -325
rect -29 -386 29 -359
rect 99 287 157 314
rect 99 253 111 287
rect 145 253 157 287
rect 99 219 157 253
rect 99 185 111 219
rect 145 185 157 219
rect 99 151 157 185
rect 99 117 111 151
rect 145 117 157 151
rect 99 83 157 117
rect 99 49 111 83
rect 145 49 157 83
rect 99 15 157 49
rect 99 -19 111 15
rect 145 -19 157 15
rect 99 -53 157 -19
rect 99 -87 111 -53
rect 145 -87 157 -53
rect 99 -121 157 -87
rect 99 -155 111 -121
rect 145 -155 157 -121
rect 99 -189 157 -155
rect 99 -223 111 -189
rect 145 -223 157 -189
rect 99 -257 157 -223
rect 99 -291 111 -257
rect 145 -291 157 -257
rect 99 -325 157 -291
rect 99 -359 111 -325
rect 145 -359 157 -325
rect 99 -386 157 -359
rect 227 287 285 314
rect 227 253 239 287
rect 273 253 285 287
rect 227 219 285 253
rect 227 185 239 219
rect 273 185 285 219
rect 227 151 285 185
rect 227 117 239 151
rect 273 117 285 151
rect 227 83 285 117
rect 227 49 239 83
rect 273 49 285 83
rect 227 15 285 49
rect 227 -19 239 15
rect 273 -19 285 15
rect 227 -53 285 -19
rect 227 -87 239 -53
rect 273 -87 285 -53
rect 227 -121 285 -87
rect 227 -155 239 -121
rect 273 -155 285 -121
rect 227 -189 285 -155
rect 227 -223 239 -189
rect 273 -223 285 -189
rect 227 -257 285 -223
rect 227 -291 239 -257
rect 273 -291 285 -257
rect 227 -325 285 -291
rect 227 -359 239 -325
rect 273 -359 285 -325
rect 227 -386 285 -359
rect 355 287 413 314
rect 355 253 367 287
rect 401 253 413 287
rect 355 219 413 253
rect 355 185 367 219
rect 401 185 413 219
rect 355 151 413 185
rect 355 117 367 151
rect 401 117 413 151
rect 355 83 413 117
rect 355 49 367 83
rect 401 49 413 83
rect 355 15 413 49
rect 355 -19 367 15
rect 401 -19 413 15
rect 355 -53 413 -19
rect 355 -87 367 -53
rect 401 -87 413 -53
rect 355 -121 413 -87
rect 355 -155 367 -121
rect 401 -155 413 -121
rect 355 -189 413 -155
rect 355 -223 367 -189
rect 401 -223 413 -189
rect 355 -257 413 -223
rect 355 -291 367 -257
rect 401 -291 413 -257
rect 355 -325 413 -291
rect 355 -359 367 -325
rect 401 -359 413 -325
rect 355 -386 413 -359
rect 483 287 541 314
rect 483 253 495 287
rect 529 253 541 287
rect 483 219 541 253
rect 483 185 495 219
rect 529 185 541 219
rect 483 151 541 185
rect 483 117 495 151
rect 529 117 541 151
rect 483 83 541 117
rect 483 49 495 83
rect 529 49 541 83
rect 483 15 541 49
rect 483 -19 495 15
rect 529 -19 541 15
rect 483 -53 541 -19
rect 483 -87 495 -53
rect 529 -87 541 -53
rect 483 -121 541 -87
rect 483 -155 495 -121
rect 529 -155 541 -121
rect 483 -189 541 -155
rect 483 -223 495 -189
rect 529 -223 541 -189
rect 483 -257 541 -223
rect 483 -291 495 -257
rect 529 -291 541 -257
rect 483 -325 541 -291
rect 483 -359 495 -325
rect 529 -359 541 -325
rect 483 -386 541 -359
rect 611 287 669 314
rect 611 253 623 287
rect 657 253 669 287
rect 611 219 669 253
rect 611 185 623 219
rect 657 185 669 219
rect 611 151 669 185
rect 611 117 623 151
rect 657 117 669 151
rect 611 83 669 117
rect 611 49 623 83
rect 657 49 669 83
rect 611 15 669 49
rect 611 -19 623 15
rect 657 -19 669 15
rect 611 -53 669 -19
rect 611 -87 623 -53
rect 657 -87 669 -53
rect 611 -121 669 -87
rect 611 -155 623 -121
rect 657 -155 669 -121
rect 611 -189 669 -155
rect 611 -223 623 -189
rect 657 -223 669 -189
rect 611 -257 669 -223
rect 611 -291 623 -257
rect 657 -291 669 -257
rect 611 -325 669 -291
rect 611 -359 623 -325
rect 657 -359 669 -325
rect 611 -386 669 -359
rect 739 287 797 314
rect 739 253 751 287
rect 785 253 797 287
rect 739 219 797 253
rect 739 185 751 219
rect 785 185 797 219
rect 739 151 797 185
rect 739 117 751 151
rect 785 117 797 151
rect 739 83 797 117
rect 739 49 751 83
rect 785 49 797 83
rect 739 15 797 49
rect 739 -19 751 15
rect 785 -19 797 15
rect 739 -53 797 -19
rect 739 -87 751 -53
rect 785 -87 797 -53
rect 739 -121 797 -87
rect 739 -155 751 -121
rect 785 -155 797 -121
rect 739 -189 797 -155
rect 739 -223 751 -189
rect 785 -223 797 -189
rect 739 -257 797 -223
rect 739 -291 751 -257
rect 785 -291 797 -257
rect 739 -325 797 -291
rect 739 -359 751 -325
rect 785 -359 797 -325
rect 739 -386 797 -359
rect 867 287 925 314
rect 867 253 879 287
rect 913 253 925 287
rect 867 219 925 253
rect 867 185 879 219
rect 913 185 925 219
rect 867 151 925 185
rect 867 117 879 151
rect 913 117 925 151
rect 867 83 925 117
rect 867 49 879 83
rect 913 49 925 83
rect 867 15 925 49
rect 867 -19 879 15
rect 913 -19 925 15
rect 867 -53 925 -19
rect 867 -87 879 -53
rect 913 -87 925 -53
rect 867 -121 925 -87
rect 867 -155 879 -121
rect 913 -155 925 -121
rect 867 -189 925 -155
rect 867 -223 879 -189
rect 913 -223 925 -189
rect 867 -257 925 -223
rect 867 -291 879 -257
rect 913 -291 925 -257
rect 867 -325 925 -291
rect 867 -359 879 -325
rect 913 -359 925 -325
rect 867 -386 925 -359
rect 995 287 1053 314
rect 995 253 1007 287
rect 1041 253 1053 287
rect 995 219 1053 253
rect 995 185 1007 219
rect 1041 185 1053 219
rect 995 151 1053 185
rect 995 117 1007 151
rect 1041 117 1053 151
rect 995 83 1053 117
rect 995 49 1007 83
rect 1041 49 1053 83
rect 995 15 1053 49
rect 995 -19 1007 15
rect 1041 -19 1053 15
rect 995 -53 1053 -19
rect 995 -87 1007 -53
rect 1041 -87 1053 -53
rect 995 -121 1053 -87
rect 995 -155 1007 -121
rect 1041 -155 1053 -121
rect 995 -189 1053 -155
rect 995 -223 1007 -189
rect 1041 -223 1053 -189
rect 995 -257 1053 -223
rect 995 -291 1007 -257
rect 1041 -291 1053 -257
rect 995 -325 1053 -291
rect 995 -359 1007 -325
rect 1041 -359 1053 -325
rect 995 -386 1053 -359
rect 1123 287 1181 314
rect 1123 253 1135 287
rect 1169 253 1181 287
rect 1123 219 1181 253
rect 1123 185 1135 219
rect 1169 185 1181 219
rect 1123 151 1181 185
rect 1123 117 1135 151
rect 1169 117 1181 151
rect 1123 83 1181 117
rect 1123 49 1135 83
rect 1169 49 1181 83
rect 1123 15 1181 49
rect 1123 -19 1135 15
rect 1169 -19 1181 15
rect 1123 -53 1181 -19
rect 1123 -87 1135 -53
rect 1169 -87 1181 -53
rect 1123 -121 1181 -87
rect 1123 -155 1135 -121
rect 1169 -155 1181 -121
rect 1123 -189 1181 -155
rect 1123 -223 1135 -189
rect 1169 -223 1181 -189
rect 1123 -257 1181 -223
rect 1123 -291 1135 -257
rect 1169 -291 1181 -257
rect 1123 -325 1181 -291
rect 1123 -359 1135 -325
rect 1169 -359 1181 -325
rect 1123 -386 1181 -359
rect 1251 287 1309 314
rect 1251 253 1263 287
rect 1297 253 1309 287
rect 1251 219 1309 253
rect 1251 185 1263 219
rect 1297 185 1309 219
rect 1251 151 1309 185
rect 1251 117 1263 151
rect 1297 117 1309 151
rect 1251 83 1309 117
rect 1251 49 1263 83
rect 1297 49 1309 83
rect 1251 15 1309 49
rect 1251 -19 1263 15
rect 1297 -19 1309 15
rect 1251 -53 1309 -19
rect 1251 -87 1263 -53
rect 1297 -87 1309 -53
rect 1251 -121 1309 -87
rect 1251 -155 1263 -121
rect 1297 -155 1309 -121
rect 1251 -189 1309 -155
rect 1251 -223 1263 -189
rect 1297 -223 1309 -189
rect 1251 -257 1309 -223
rect 1251 -291 1263 -257
rect 1297 -291 1309 -257
rect 1251 -325 1309 -291
rect 1251 -359 1263 -325
rect 1297 -359 1309 -325
rect 1251 -386 1309 -359
rect 1379 287 1437 314
rect 1379 253 1391 287
rect 1425 253 1437 287
rect 1379 219 1437 253
rect 1379 185 1391 219
rect 1425 185 1437 219
rect 1379 151 1437 185
rect 1379 117 1391 151
rect 1425 117 1437 151
rect 1379 83 1437 117
rect 1379 49 1391 83
rect 1425 49 1437 83
rect 1379 15 1437 49
rect 1379 -19 1391 15
rect 1425 -19 1437 15
rect 1379 -53 1437 -19
rect 1379 -87 1391 -53
rect 1425 -87 1437 -53
rect 1379 -121 1437 -87
rect 1379 -155 1391 -121
rect 1425 -155 1437 -121
rect 1379 -189 1437 -155
rect 1379 -223 1391 -189
rect 1425 -223 1437 -189
rect 1379 -257 1437 -223
rect 1379 -291 1391 -257
rect 1425 -291 1437 -257
rect 1379 -325 1437 -291
rect 1379 -359 1391 -325
rect 1425 -359 1437 -325
rect 1379 -386 1437 -359
rect 1507 287 1565 314
rect 1507 253 1519 287
rect 1553 253 1565 287
rect 1507 219 1565 253
rect 1507 185 1519 219
rect 1553 185 1565 219
rect 1507 151 1565 185
rect 1507 117 1519 151
rect 1553 117 1565 151
rect 1507 83 1565 117
rect 1507 49 1519 83
rect 1553 49 1565 83
rect 1507 15 1565 49
rect 1507 -19 1519 15
rect 1553 -19 1565 15
rect 1507 -53 1565 -19
rect 1507 -87 1519 -53
rect 1553 -87 1565 -53
rect 1507 -121 1565 -87
rect 1507 -155 1519 -121
rect 1553 -155 1565 -121
rect 1507 -189 1565 -155
rect 1507 -223 1519 -189
rect 1553 -223 1565 -189
rect 1507 -257 1565 -223
rect 1507 -291 1519 -257
rect 1553 -291 1565 -257
rect 1507 -325 1565 -291
rect 1507 -359 1519 -325
rect 1553 -359 1565 -325
rect 1507 -386 1565 -359
rect 1635 287 1693 314
rect 1635 253 1647 287
rect 1681 253 1693 287
rect 1635 219 1693 253
rect 1635 185 1647 219
rect 1681 185 1693 219
rect 1635 151 1693 185
rect 1635 117 1647 151
rect 1681 117 1693 151
rect 1635 83 1693 117
rect 1635 49 1647 83
rect 1681 49 1693 83
rect 1635 15 1693 49
rect 1635 -19 1647 15
rect 1681 -19 1693 15
rect 1635 -53 1693 -19
rect 1635 -87 1647 -53
rect 1681 -87 1693 -53
rect 1635 -121 1693 -87
rect 1635 -155 1647 -121
rect 1681 -155 1693 -121
rect 1635 -189 1693 -155
rect 1635 -223 1647 -189
rect 1681 -223 1693 -189
rect 1635 -257 1693 -223
rect 1635 -291 1647 -257
rect 1681 -291 1693 -257
rect 1635 -325 1693 -291
rect 1635 -359 1647 -325
rect 1681 -359 1693 -325
rect 1635 -386 1693 -359
rect 1763 287 1821 314
rect 1763 253 1775 287
rect 1809 253 1821 287
rect 1763 219 1821 253
rect 1763 185 1775 219
rect 1809 185 1821 219
rect 1763 151 1821 185
rect 1763 117 1775 151
rect 1809 117 1821 151
rect 1763 83 1821 117
rect 1763 49 1775 83
rect 1809 49 1821 83
rect 1763 15 1821 49
rect 1763 -19 1775 15
rect 1809 -19 1821 15
rect 1763 -53 1821 -19
rect 1763 -87 1775 -53
rect 1809 -87 1821 -53
rect 1763 -121 1821 -87
rect 1763 -155 1775 -121
rect 1809 -155 1821 -121
rect 1763 -189 1821 -155
rect 1763 -223 1775 -189
rect 1809 -223 1821 -189
rect 1763 -257 1821 -223
rect 1763 -291 1775 -257
rect 1809 -291 1821 -257
rect 1763 -325 1821 -291
rect 1763 -359 1775 -325
rect 1809 -359 1821 -325
rect 1763 -386 1821 -359
rect 1891 287 1949 314
rect 1891 253 1903 287
rect 1937 253 1949 287
rect 1891 219 1949 253
rect 1891 185 1903 219
rect 1937 185 1949 219
rect 1891 151 1949 185
rect 1891 117 1903 151
rect 1937 117 1949 151
rect 1891 83 1949 117
rect 1891 49 1903 83
rect 1937 49 1949 83
rect 1891 15 1949 49
rect 1891 -19 1903 15
rect 1937 -19 1949 15
rect 1891 -53 1949 -19
rect 1891 -87 1903 -53
rect 1937 -87 1949 -53
rect 1891 -121 1949 -87
rect 1891 -155 1903 -121
rect 1937 -155 1949 -121
rect 1891 -189 1949 -155
rect 1891 -223 1903 -189
rect 1937 -223 1949 -189
rect 1891 -257 1949 -223
rect 1891 -291 1903 -257
rect 1937 -291 1949 -257
rect 1891 -325 1949 -291
rect 1891 -359 1903 -325
rect 1937 -359 1949 -325
rect 1891 -386 1949 -359
rect 2019 287 2077 314
rect 2019 253 2031 287
rect 2065 253 2077 287
rect 2019 219 2077 253
rect 2019 185 2031 219
rect 2065 185 2077 219
rect 2019 151 2077 185
rect 2019 117 2031 151
rect 2065 117 2077 151
rect 2019 83 2077 117
rect 2019 49 2031 83
rect 2065 49 2077 83
rect 2019 15 2077 49
rect 2019 -19 2031 15
rect 2065 -19 2077 15
rect 2019 -53 2077 -19
rect 2019 -87 2031 -53
rect 2065 -87 2077 -53
rect 2019 -121 2077 -87
rect 2019 -155 2031 -121
rect 2065 -155 2077 -121
rect 2019 -189 2077 -155
rect 2019 -223 2031 -189
rect 2065 -223 2077 -189
rect 2019 -257 2077 -223
rect 2019 -291 2031 -257
rect 2065 -291 2077 -257
rect 2019 -325 2077 -291
rect 2019 -359 2031 -325
rect 2065 -359 2077 -325
rect 2019 -386 2077 -359
rect 2147 287 2205 314
rect 2147 253 2159 287
rect 2193 253 2205 287
rect 2147 219 2205 253
rect 2147 185 2159 219
rect 2193 185 2205 219
rect 2147 151 2205 185
rect 2147 117 2159 151
rect 2193 117 2205 151
rect 2147 83 2205 117
rect 2147 49 2159 83
rect 2193 49 2205 83
rect 2147 15 2205 49
rect 2147 -19 2159 15
rect 2193 -19 2205 15
rect 2147 -53 2205 -19
rect 2147 -87 2159 -53
rect 2193 -87 2205 -53
rect 2147 -121 2205 -87
rect 2147 -155 2159 -121
rect 2193 -155 2205 -121
rect 2147 -189 2205 -155
rect 2147 -223 2159 -189
rect 2193 -223 2205 -189
rect 2147 -257 2205 -223
rect 2147 -291 2159 -257
rect 2193 -291 2205 -257
rect 2147 -325 2205 -291
rect 2147 -359 2159 -325
rect 2193 -359 2205 -325
rect 2147 -386 2205 -359
rect 2275 287 2333 314
rect 2275 253 2287 287
rect 2321 253 2333 287
rect 2275 219 2333 253
rect 2275 185 2287 219
rect 2321 185 2333 219
rect 2275 151 2333 185
rect 2275 117 2287 151
rect 2321 117 2333 151
rect 2275 83 2333 117
rect 2275 49 2287 83
rect 2321 49 2333 83
rect 2275 15 2333 49
rect 2275 -19 2287 15
rect 2321 -19 2333 15
rect 2275 -53 2333 -19
rect 2275 -87 2287 -53
rect 2321 -87 2333 -53
rect 2275 -121 2333 -87
rect 2275 -155 2287 -121
rect 2321 -155 2333 -121
rect 2275 -189 2333 -155
rect 2275 -223 2287 -189
rect 2321 -223 2333 -189
rect 2275 -257 2333 -223
rect 2275 -291 2287 -257
rect 2321 -291 2333 -257
rect 2275 -325 2333 -291
rect 2275 -359 2287 -325
rect 2321 -359 2333 -325
rect 2275 -386 2333 -359
rect 2403 287 2461 314
rect 2403 253 2415 287
rect 2449 253 2461 287
rect 2403 219 2461 253
rect 2403 185 2415 219
rect 2449 185 2461 219
rect 2403 151 2461 185
rect 2403 117 2415 151
rect 2449 117 2461 151
rect 2403 83 2461 117
rect 2403 49 2415 83
rect 2449 49 2461 83
rect 2403 15 2461 49
rect 2403 -19 2415 15
rect 2449 -19 2461 15
rect 2403 -53 2461 -19
rect 2403 -87 2415 -53
rect 2449 -87 2461 -53
rect 2403 -121 2461 -87
rect 2403 -155 2415 -121
rect 2449 -155 2461 -121
rect 2403 -189 2461 -155
rect 2403 -223 2415 -189
rect 2449 -223 2461 -189
rect 2403 -257 2461 -223
rect 2403 -291 2415 -257
rect 2449 -291 2461 -257
rect 2403 -325 2461 -291
rect 2403 -359 2415 -325
rect 2449 -359 2461 -325
rect 2403 -386 2461 -359
rect 2531 287 2589 314
rect 2531 253 2543 287
rect 2577 253 2589 287
rect 2531 219 2589 253
rect 2531 185 2543 219
rect 2577 185 2589 219
rect 2531 151 2589 185
rect 2531 117 2543 151
rect 2577 117 2589 151
rect 2531 83 2589 117
rect 2531 49 2543 83
rect 2577 49 2589 83
rect 2531 15 2589 49
rect 2531 -19 2543 15
rect 2577 -19 2589 15
rect 2531 -53 2589 -19
rect 2531 -87 2543 -53
rect 2577 -87 2589 -53
rect 2531 -121 2589 -87
rect 2531 -155 2543 -121
rect 2577 -155 2589 -121
rect 2531 -189 2589 -155
rect 2531 -223 2543 -189
rect 2577 -223 2589 -189
rect 2531 -257 2589 -223
rect 2531 -291 2543 -257
rect 2577 -291 2589 -257
rect 2531 -325 2589 -291
rect 2531 -359 2543 -325
rect 2577 -359 2589 -325
rect 2531 -386 2589 -359
<< pdiffc >>
rect -2577 253 -2543 287
rect -2577 185 -2543 219
rect -2577 117 -2543 151
rect -2577 49 -2543 83
rect -2577 -19 -2543 15
rect -2577 -87 -2543 -53
rect -2577 -155 -2543 -121
rect -2577 -223 -2543 -189
rect -2577 -291 -2543 -257
rect -2577 -359 -2543 -325
rect -2449 253 -2415 287
rect -2449 185 -2415 219
rect -2449 117 -2415 151
rect -2449 49 -2415 83
rect -2449 -19 -2415 15
rect -2449 -87 -2415 -53
rect -2449 -155 -2415 -121
rect -2449 -223 -2415 -189
rect -2449 -291 -2415 -257
rect -2449 -359 -2415 -325
rect -2321 253 -2287 287
rect -2321 185 -2287 219
rect -2321 117 -2287 151
rect -2321 49 -2287 83
rect -2321 -19 -2287 15
rect -2321 -87 -2287 -53
rect -2321 -155 -2287 -121
rect -2321 -223 -2287 -189
rect -2321 -291 -2287 -257
rect -2321 -359 -2287 -325
rect -2193 253 -2159 287
rect -2193 185 -2159 219
rect -2193 117 -2159 151
rect -2193 49 -2159 83
rect -2193 -19 -2159 15
rect -2193 -87 -2159 -53
rect -2193 -155 -2159 -121
rect -2193 -223 -2159 -189
rect -2193 -291 -2159 -257
rect -2193 -359 -2159 -325
rect -2065 253 -2031 287
rect -2065 185 -2031 219
rect -2065 117 -2031 151
rect -2065 49 -2031 83
rect -2065 -19 -2031 15
rect -2065 -87 -2031 -53
rect -2065 -155 -2031 -121
rect -2065 -223 -2031 -189
rect -2065 -291 -2031 -257
rect -2065 -359 -2031 -325
rect -1937 253 -1903 287
rect -1937 185 -1903 219
rect -1937 117 -1903 151
rect -1937 49 -1903 83
rect -1937 -19 -1903 15
rect -1937 -87 -1903 -53
rect -1937 -155 -1903 -121
rect -1937 -223 -1903 -189
rect -1937 -291 -1903 -257
rect -1937 -359 -1903 -325
rect -1809 253 -1775 287
rect -1809 185 -1775 219
rect -1809 117 -1775 151
rect -1809 49 -1775 83
rect -1809 -19 -1775 15
rect -1809 -87 -1775 -53
rect -1809 -155 -1775 -121
rect -1809 -223 -1775 -189
rect -1809 -291 -1775 -257
rect -1809 -359 -1775 -325
rect -1681 253 -1647 287
rect -1681 185 -1647 219
rect -1681 117 -1647 151
rect -1681 49 -1647 83
rect -1681 -19 -1647 15
rect -1681 -87 -1647 -53
rect -1681 -155 -1647 -121
rect -1681 -223 -1647 -189
rect -1681 -291 -1647 -257
rect -1681 -359 -1647 -325
rect -1553 253 -1519 287
rect -1553 185 -1519 219
rect -1553 117 -1519 151
rect -1553 49 -1519 83
rect -1553 -19 -1519 15
rect -1553 -87 -1519 -53
rect -1553 -155 -1519 -121
rect -1553 -223 -1519 -189
rect -1553 -291 -1519 -257
rect -1553 -359 -1519 -325
rect -1425 253 -1391 287
rect -1425 185 -1391 219
rect -1425 117 -1391 151
rect -1425 49 -1391 83
rect -1425 -19 -1391 15
rect -1425 -87 -1391 -53
rect -1425 -155 -1391 -121
rect -1425 -223 -1391 -189
rect -1425 -291 -1391 -257
rect -1425 -359 -1391 -325
rect -1297 253 -1263 287
rect -1297 185 -1263 219
rect -1297 117 -1263 151
rect -1297 49 -1263 83
rect -1297 -19 -1263 15
rect -1297 -87 -1263 -53
rect -1297 -155 -1263 -121
rect -1297 -223 -1263 -189
rect -1297 -291 -1263 -257
rect -1297 -359 -1263 -325
rect -1169 253 -1135 287
rect -1169 185 -1135 219
rect -1169 117 -1135 151
rect -1169 49 -1135 83
rect -1169 -19 -1135 15
rect -1169 -87 -1135 -53
rect -1169 -155 -1135 -121
rect -1169 -223 -1135 -189
rect -1169 -291 -1135 -257
rect -1169 -359 -1135 -325
rect -1041 253 -1007 287
rect -1041 185 -1007 219
rect -1041 117 -1007 151
rect -1041 49 -1007 83
rect -1041 -19 -1007 15
rect -1041 -87 -1007 -53
rect -1041 -155 -1007 -121
rect -1041 -223 -1007 -189
rect -1041 -291 -1007 -257
rect -1041 -359 -1007 -325
rect -913 253 -879 287
rect -913 185 -879 219
rect -913 117 -879 151
rect -913 49 -879 83
rect -913 -19 -879 15
rect -913 -87 -879 -53
rect -913 -155 -879 -121
rect -913 -223 -879 -189
rect -913 -291 -879 -257
rect -913 -359 -879 -325
rect -785 253 -751 287
rect -785 185 -751 219
rect -785 117 -751 151
rect -785 49 -751 83
rect -785 -19 -751 15
rect -785 -87 -751 -53
rect -785 -155 -751 -121
rect -785 -223 -751 -189
rect -785 -291 -751 -257
rect -785 -359 -751 -325
rect -657 253 -623 287
rect -657 185 -623 219
rect -657 117 -623 151
rect -657 49 -623 83
rect -657 -19 -623 15
rect -657 -87 -623 -53
rect -657 -155 -623 -121
rect -657 -223 -623 -189
rect -657 -291 -623 -257
rect -657 -359 -623 -325
rect -529 253 -495 287
rect -529 185 -495 219
rect -529 117 -495 151
rect -529 49 -495 83
rect -529 -19 -495 15
rect -529 -87 -495 -53
rect -529 -155 -495 -121
rect -529 -223 -495 -189
rect -529 -291 -495 -257
rect -529 -359 -495 -325
rect -401 253 -367 287
rect -401 185 -367 219
rect -401 117 -367 151
rect -401 49 -367 83
rect -401 -19 -367 15
rect -401 -87 -367 -53
rect -401 -155 -367 -121
rect -401 -223 -367 -189
rect -401 -291 -367 -257
rect -401 -359 -367 -325
rect -273 253 -239 287
rect -273 185 -239 219
rect -273 117 -239 151
rect -273 49 -239 83
rect -273 -19 -239 15
rect -273 -87 -239 -53
rect -273 -155 -239 -121
rect -273 -223 -239 -189
rect -273 -291 -239 -257
rect -273 -359 -239 -325
rect -145 253 -111 287
rect -145 185 -111 219
rect -145 117 -111 151
rect -145 49 -111 83
rect -145 -19 -111 15
rect -145 -87 -111 -53
rect -145 -155 -111 -121
rect -145 -223 -111 -189
rect -145 -291 -111 -257
rect -145 -359 -111 -325
rect -17 253 17 287
rect -17 185 17 219
rect -17 117 17 151
rect -17 49 17 83
rect -17 -19 17 15
rect -17 -87 17 -53
rect -17 -155 17 -121
rect -17 -223 17 -189
rect -17 -291 17 -257
rect -17 -359 17 -325
rect 111 253 145 287
rect 111 185 145 219
rect 111 117 145 151
rect 111 49 145 83
rect 111 -19 145 15
rect 111 -87 145 -53
rect 111 -155 145 -121
rect 111 -223 145 -189
rect 111 -291 145 -257
rect 111 -359 145 -325
rect 239 253 273 287
rect 239 185 273 219
rect 239 117 273 151
rect 239 49 273 83
rect 239 -19 273 15
rect 239 -87 273 -53
rect 239 -155 273 -121
rect 239 -223 273 -189
rect 239 -291 273 -257
rect 239 -359 273 -325
rect 367 253 401 287
rect 367 185 401 219
rect 367 117 401 151
rect 367 49 401 83
rect 367 -19 401 15
rect 367 -87 401 -53
rect 367 -155 401 -121
rect 367 -223 401 -189
rect 367 -291 401 -257
rect 367 -359 401 -325
rect 495 253 529 287
rect 495 185 529 219
rect 495 117 529 151
rect 495 49 529 83
rect 495 -19 529 15
rect 495 -87 529 -53
rect 495 -155 529 -121
rect 495 -223 529 -189
rect 495 -291 529 -257
rect 495 -359 529 -325
rect 623 253 657 287
rect 623 185 657 219
rect 623 117 657 151
rect 623 49 657 83
rect 623 -19 657 15
rect 623 -87 657 -53
rect 623 -155 657 -121
rect 623 -223 657 -189
rect 623 -291 657 -257
rect 623 -359 657 -325
rect 751 253 785 287
rect 751 185 785 219
rect 751 117 785 151
rect 751 49 785 83
rect 751 -19 785 15
rect 751 -87 785 -53
rect 751 -155 785 -121
rect 751 -223 785 -189
rect 751 -291 785 -257
rect 751 -359 785 -325
rect 879 253 913 287
rect 879 185 913 219
rect 879 117 913 151
rect 879 49 913 83
rect 879 -19 913 15
rect 879 -87 913 -53
rect 879 -155 913 -121
rect 879 -223 913 -189
rect 879 -291 913 -257
rect 879 -359 913 -325
rect 1007 253 1041 287
rect 1007 185 1041 219
rect 1007 117 1041 151
rect 1007 49 1041 83
rect 1007 -19 1041 15
rect 1007 -87 1041 -53
rect 1007 -155 1041 -121
rect 1007 -223 1041 -189
rect 1007 -291 1041 -257
rect 1007 -359 1041 -325
rect 1135 253 1169 287
rect 1135 185 1169 219
rect 1135 117 1169 151
rect 1135 49 1169 83
rect 1135 -19 1169 15
rect 1135 -87 1169 -53
rect 1135 -155 1169 -121
rect 1135 -223 1169 -189
rect 1135 -291 1169 -257
rect 1135 -359 1169 -325
rect 1263 253 1297 287
rect 1263 185 1297 219
rect 1263 117 1297 151
rect 1263 49 1297 83
rect 1263 -19 1297 15
rect 1263 -87 1297 -53
rect 1263 -155 1297 -121
rect 1263 -223 1297 -189
rect 1263 -291 1297 -257
rect 1263 -359 1297 -325
rect 1391 253 1425 287
rect 1391 185 1425 219
rect 1391 117 1425 151
rect 1391 49 1425 83
rect 1391 -19 1425 15
rect 1391 -87 1425 -53
rect 1391 -155 1425 -121
rect 1391 -223 1425 -189
rect 1391 -291 1425 -257
rect 1391 -359 1425 -325
rect 1519 253 1553 287
rect 1519 185 1553 219
rect 1519 117 1553 151
rect 1519 49 1553 83
rect 1519 -19 1553 15
rect 1519 -87 1553 -53
rect 1519 -155 1553 -121
rect 1519 -223 1553 -189
rect 1519 -291 1553 -257
rect 1519 -359 1553 -325
rect 1647 253 1681 287
rect 1647 185 1681 219
rect 1647 117 1681 151
rect 1647 49 1681 83
rect 1647 -19 1681 15
rect 1647 -87 1681 -53
rect 1647 -155 1681 -121
rect 1647 -223 1681 -189
rect 1647 -291 1681 -257
rect 1647 -359 1681 -325
rect 1775 253 1809 287
rect 1775 185 1809 219
rect 1775 117 1809 151
rect 1775 49 1809 83
rect 1775 -19 1809 15
rect 1775 -87 1809 -53
rect 1775 -155 1809 -121
rect 1775 -223 1809 -189
rect 1775 -291 1809 -257
rect 1775 -359 1809 -325
rect 1903 253 1937 287
rect 1903 185 1937 219
rect 1903 117 1937 151
rect 1903 49 1937 83
rect 1903 -19 1937 15
rect 1903 -87 1937 -53
rect 1903 -155 1937 -121
rect 1903 -223 1937 -189
rect 1903 -291 1937 -257
rect 1903 -359 1937 -325
rect 2031 253 2065 287
rect 2031 185 2065 219
rect 2031 117 2065 151
rect 2031 49 2065 83
rect 2031 -19 2065 15
rect 2031 -87 2065 -53
rect 2031 -155 2065 -121
rect 2031 -223 2065 -189
rect 2031 -291 2065 -257
rect 2031 -359 2065 -325
rect 2159 253 2193 287
rect 2159 185 2193 219
rect 2159 117 2193 151
rect 2159 49 2193 83
rect 2159 -19 2193 15
rect 2159 -87 2193 -53
rect 2159 -155 2193 -121
rect 2159 -223 2193 -189
rect 2159 -291 2193 -257
rect 2159 -359 2193 -325
rect 2287 253 2321 287
rect 2287 185 2321 219
rect 2287 117 2321 151
rect 2287 49 2321 83
rect 2287 -19 2321 15
rect 2287 -87 2321 -53
rect 2287 -155 2321 -121
rect 2287 -223 2321 -189
rect 2287 -291 2321 -257
rect 2287 -359 2321 -325
rect 2415 253 2449 287
rect 2415 185 2449 219
rect 2415 117 2449 151
rect 2415 49 2449 83
rect 2415 -19 2449 15
rect 2415 -87 2449 -53
rect 2415 -155 2449 -121
rect 2415 -223 2449 -189
rect 2415 -291 2449 -257
rect 2415 -359 2449 -325
rect 2543 253 2577 287
rect 2543 185 2577 219
rect 2543 117 2577 151
rect 2543 49 2577 83
rect 2543 -19 2577 15
rect 2543 -87 2577 -53
rect 2543 -155 2577 -121
rect 2543 -223 2577 -189
rect 2543 -291 2577 -257
rect 2543 -359 2577 -325
<< nsubdiff >>
rect -2691 464 -2567 498
rect -2533 464 -2499 498
rect -2465 464 -2431 498
rect -2397 464 -2363 498
rect -2329 464 -2295 498
rect -2261 464 -2227 498
rect -2193 464 -2159 498
rect -2125 464 -2091 498
rect -2057 464 -2023 498
rect -1989 464 -1955 498
rect -1921 464 -1887 498
rect -1853 464 -1819 498
rect -1785 464 -1751 498
rect -1717 464 -1683 498
rect -1649 464 -1615 498
rect -1581 464 -1547 498
rect -1513 464 -1479 498
rect -1445 464 -1411 498
rect -1377 464 -1343 498
rect -1309 464 -1275 498
rect -1241 464 -1207 498
rect -1173 464 -1139 498
rect -1105 464 -1071 498
rect -1037 464 -1003 498
rect -969 464 -935 498
rect -901 464 -867 498
rect -833 464 -799 498
rect -765 464 -731 498
rect -697 464 -663 498
rect -629 464 -595 498
rect -561 464 -527 498
rect -493 464 -459 498
rect -425 464 -391 498
rect -357 464 -323 498
rect -289 464 -255 498
rect -221 464 -187 498
rect -153 464 -119 498
rect -85 464 -51 498
rect -17 464 17 498
rect 51 464 85 498
rect 119 464 153 498
rect 187 464 221 498
rect 255 464 289 498
rect 323 464 357 498
rect 391 464 425 498
rect 459 464 493 498
rect 527 464 561 498
rect 595 464 629 498
rect 663 464 697 498
rect 731 464 765 498
rect 799 464 833 498
rect 867 464 901 498
rect 935 464 969 498
rect 1003 464 1037 498
rect 1071 464 1105 498
rect 1139 464 1173 498
rect 1207 464 1241 498
rect 1275 464 1309 498
rect 1343 464 1377 498
rect 1411 464 1445 498
rect 1479 464 1513 498
rect 1547 464 1581 498
rect 1615 464 1649 498
rect 1683 464 1717 498
rect 1751 464 1785 498
rect 1819 464 1853 498
rect 1887 464 1921 498
rect 1955 464 1989 498
rect 2023 464 2057 498
rect 2091 464 2125 498
rect 2159 464 2193 498
rect 2227 464 2261 498
rect 2295 464 2329 498
rect 2363 464 2397 498
rect 2431 464 2465 498
rect 2499 464 2533 498
rect 2567 464 2691 498
rect -2691 391 -2657 464
rect -2691 323 -2657 357
rect 2657 391 2691 464
rect 2657 323 2691 357
rect -2691 255 -2657 289
rect -2691 187 -2657 221
rect -2691 119 -2657 153
rect -2691 51 -2657 85
rect -2691 -17 -2657 17
rect -2691 -85 -2657 -51
rect -2691 -153 -2657 -119
rect -2691 -221 -2657 -187
rect -2691 -289 -2657 -255
rect -2691 -357 -2657 -323
rect 2657 255 2691 289
rect 2657 187 2691 221
rect 2657 119 2691 153
rect 2657 51 2691 85
rect 2657 -17 2691 17
rect 2657 -85 2691 -51
rect 2657 -153 2691 -119
rect 2657 -221 2691 -187
rect 2657 -289 2691 -255
rect 2657 -357 2691 -323
rect -2691 -464 -2657 -391
rect 2657 -464 2691 -391
rect -2691 -498 -2567 -464
rect -2533 -498 -2499 -464
rect -2465 -498 -2431 -464
rect -2397 -498 -2363 -464
rect -2329 -498 -2295 -464
rect -2261 -498 -2227 -464
rect -2193 -498 -2159 -464
rect -2125 -498 -2091 -464
rect -2057 -498 -2023 -464
rect -1989 -498 -1955 -464
rect -1921 -498 -1887 -464
rect -1853 -498 -1819 -464
rect -1785 -498 -1751 -464
rect -1717 -498 -1683 -464
rect -1649 -498 -1615 -464
rect -1581 -498 -1547 -464
rect -1513 -498 -1479 -464
rect -1445 -498 -1411 -464
rect -1377 -498 -1343 -464
rect -1309 -498 -1275 -464
rect -1241 -498 -1207 -464
rect -1173 -498 -1139 -464
rect -1105 -498 -1071 -464
rect -1037 -498 -1003 -464
rect -969 -498 -935 -464
rect -901 -498 -867 -464
rect -833 -498 -799 -464
rect -765 -498 -731 -464
rect -697 -498 -663 -464
rect -629 -498 -595 -464
rect -561 -498 -527 -464
rect -493 -498 -459 -464
rect -425 -498 -391 -464
rect -357 -498 -323 -464
rect -289 -498 -255 -464
rect -221 -498 -187 -464
rect -153 -498 -119 -464
rect -85 -498 -51 -464
rect -17 -498 17 -464
rect 51 -498 85 -464
rect 119 -498 153 -464
rect 187 -498 221 -464
rect 255 -498 289 -464
rect 323 -498 357 -464
rect 391 -498 425 -464
rect 459 -498 493 -464
rect 527 -498 561 -464
rect 595 -498 629 -464
rect 663 -498 697 -464
rect 731 -498 765 -464
rect 799 -498 833 -464
rect 867 -498 901 -464
rect 935 -498 969 -464
rect 1003 -498 1037 -464
rect 1071 -498 1105 -464
rect 1139 -498 1173 -464
rect 1207 -498 1241 -464
rect 1275 -498 1309 -464
rect 1343 -498 1377 -464
rect 1411 -498 1445 -464
rect 1479 -498 1513 -464
rect 1547 -498 1581 -464
rect 1615 -498 1649 -464
rect 1683 -498 1717 -464
rect 1751 -498 1785 -464
rect 1819 -498 1853 -464
rect 1887 -498 1921 -464
rect 1955 -498 1989 -464
rect 2023 -498 2057 -464
rect 2091 -498 2125 -464
rect 2159 -498 2193 -464
rect 2227 -498 2261 -464
rect 2295 -498 2329 -464
rect 2363 -498 2397 -464
rect 2431 -498 2465 -464
rect 2499 -498 2533 -464
rect 2567 -498 2691 -464
<< nsubdiffcont >>
rect -2567 464 -2533 498
rect -2499 464 -2465 498
rect -2431 464 -2397 498
rect -2363 464 -2329 498
rect -2295 464 -2261 498
rect -2227 464 -2193 498
rect -2159 464 -2125 498
rect -2091 464 -2057 498
rect -2023 464 -1989 498
rect -1955 464 -1921 498
rect -1887 464 -1853 498
rect -1819 464 -1785 498
rect -1751 464 -1717 498
rect -1683 464 -1649 498
rect -1615 464 -1581 498
rect -1547 464 -1513 498
rect -1479 464 -1445 498
rect -1411 464 -1377 498
rect -1343 464 -1309 498
rect -1275 464 -1241 498
rect -1207 464 -1173 498
rect -1139 464 -1105 498
rect -1071 464 -1037 498
rect -1003 464 -969 498
rect -935 464 -901 498
rect -867 464 -833 498
rect -799 464 -765 498
rect -731 464 -697 498
rect -663 464 -629 498
rect -595 464 -561 498
rect -527 464 -493 498
rect -459 464 -425 498
rect -391 464 -357 498
rect -323 464 -289 498
rect -255 464 -221 498
rect -187 464 -153 498
rect -119 464 -85 498
rect -51 464 -17 498
rect 17 464 51 498
rect 85 464 119 498
rect 153 464 187 498
rect 221 464 255 498
rect 289 464 323 498
rect 357 464 391 498
rect 425 464 459 498
rect 493 464 527 498
rect 561 464 595 498
rect 629 464 663 498
rect 697 464 731 498
rect 765 464 799 498
rect 833 464 867 498
rect 901 464 935 498
rect 969 464 1003 498
rect 1037 464 1071 498
rect 1105 464 1139 498
rect 1173 464 1207 498
rect 1241 464 1275 498
rect 1309 464 1343 498
rect 1377 464 1411 498
rect 1445 464 1479 498
rect 1513 464 1547 498
rect 1581 464 1615 498
rect 1649 464 1683 498
rect 1717 464 1751 498
rect 1785 464 1819 498
rect 1853 464 1887 498
rect 1921 464 1955 498
rect 1989 464 2023 498
rect 2057 464 2091 498
rect 2125 464 2159 498
rect 2193 464 2227 498
rect 2261 464 2295 498
rect 2329 464 2363 498
rect 2397 464 2431 498
rect 2465 464 2499 498
rect 2533 464 2567 498
rect -2691 357 -2657 391
rect -2691 289 -2657 323
rect 2657 357 2691 391
rect -2691 221 -2657 255
rect -2691 153 -2657 187
rect -2691 85 -2657 119
rect -2691 17 -2657 51
rect -2691 -51 -2657 -17
rect -2691 -119 -2657 -85
rect -2691 -187 -2657 -153
rect -2691 -255 -2657 -221
rect -2691 -323 -2657 -289
rect -2691 -391 -2657 -357
rect 2657 289 2691 323
rect 2657 221 2691 255
rect 2657 153 2691 187
rect 2657 85 2691 119
rect 2657 17 2691 51
rect 2657 -51 2691 -17
rect 2657 -119 2691 -85
rect 2657 -187 2691 -153
rect 2657 -255 2691 -221
rect 2657 -323 2691 -289
rect 2657 -391 2691 -357
rect -2567 -498 -2533 -464
rect -2499 -498 -2465 -464
rect -2431 -498 -2397 -464
rect -2363 -498 -2329 -464
rect -2295 -498 -2261 -464
rect -2227 -498 -2193 -464
rect -2159 -498 -2125 -464
rect -2091 -498 -2057 -464
rect -2023 -498 -1989 -464
rect -1955 -498 -1921 -464
rect -1887 -498 -1853 -464
rect -1819 -498 -1785 -464
rect -1751 -498 -1717 -464
rect -1683 -498 -1649 -464
rect -1615 -498 -1581 -464
rect -1547 -498 -1513 -464
rect -1479 -498 -1445 -464
rect -1411 -498 -1377 -464
rect -1343 -498 -1309 -464
rect -1275 -498 -1241 -464
rect -1207 -498 -1173 -464
rect -1139 -498 -1105 -464
rect -1071 -498 -1037 -464
rect -1003 -498 -969 -464
rect -935 -498 -901 -464
rect -867 -498 -833 -464
rect -799 -498 -765 -464
rect -731 -498 -697 -464
rect -663 -498 -629 -464
rect -595 -498 -561 -464
rect -527 -498 -493 -464
rect -459 -498 -425 -464
rect -391 -498 -357 -464
rect -323 -498 -289 -464
rect -255 -498 -221 -464
rect -187 -498 -153 -464
rect -119 -498 -85 -464
rect -51 -498 -17 -464
rect 17 -498 51 -464
rect 85 -498 119 -464
rect 153 -498 187 -464
rect 221 -498 255 -464
rect 289 -498 323 -464
rect 357 -498 391 -464
rect 425 -498 459 -464
rect 493 -498 527 -464
rect 561 -498 595 -464
rect 629 -498 663 -464
rect 697 -498 731 -464
rect 765 -498 799 -464
rect 833 -498 867 -464
rect 901 -498 935 -464
rect 969 -498 1003 -464
rect 1037 -498 1071 -464
rect 1105 -498 1139 -464
rect 1173 -498 1207 -464
rect 1241 -498 1275 -464
rect 1309 -498 1343 -464
rect 1377 -498 1411 -464
rect 1445 -498 1479 -464
rect 1513 -498 1547 -464
rect 1581 -498 1615 -464
rect 1649 -498 1683 -464
rect 1717 -498 1751 -464
rect 1785 -498 1819 -464
rect 1853 -498 1887 -464
rect 1921 -498 1955 -464
rect 1989 -498 2023 -464
rect 2057 -498 2091 -464
rect 2125 -498 2159 -464
rect 2193 -498 2227 -464
rect 2261 -498 2295 -464
rect 2329 -498 2363 -464
rect 2397 -498 2431 -464
rect 2465 -498 2499 -464
rect 2533 -498 2567 -464
<< poly >>
rect -2531 395 -2461 411
rect -2531 361 -2513 395
rect -2479 361 -2461 395
rect -2531 314 -2461 361
rect -2403 395 -2333 411
rect -2403 361 -2385 395
rect -2351 361 -2333 395
rect -2403 314 -2333 361
rect -2275 395 -2205 411
rect -2275 361 -2257 395
rect -2223 361 -2205 395
rect -2275 314 -2205 361
rect -2147 395 -2077 411
rect -2147 361 -2129 395
rect -2095 361 -2077 395
rect -2147 314 -2077 361
rect -2019 395 -1949 411
rect -2019 361 -2001 395
rect -1967 361 -1949 395
rect -2019 314 -1949 361
rect -1891 395 -1821 411
rect -1891 361 -1873 395
rect -1839 361 -1821 395
rect -1891 314 -1821 361
rect -1763 395 -1693 411
rect -1763 361 -1745 395
rect -1711 361 -1693 395
rect -1763 314 -1693 361
rect -1635 395 -1565 411
rect -1635 361 -1617 395
rect -1583 361 -1565 395
rect -1635 314 -1565 361
rect -1507 395 -1437 411
rect -1507 361 -1489 395
rect -1455 361 -1437 395
rect -1507 314 -1437 361
rect -1379 395 -1309 411
rect -1379 361 -1361 395
rect -1327 361 -1309 395
rect -1379 314 -1309 361
rect -1251 395 -1181 411
rect -1251 361 -1233 395
rect -1199 361 -1181 395
rect -1251 314 -1181 361
rect -1123 395 -1053 411
rect -1123 361 -1105 395
rect -1071 361 -1053 395
rect -1123 314 -1053 361
rect -995 395 -925 411
rect -995 361 -977 395
rect -943 361 -925 395
rect -995 314 -925 361
rect -867 395 -797 411
rect -867 361 -849 395
rect -815 361 -797 395
rect -867 314 -797 361
rect -739 395 -669 411
rect -739 361 -721 395
rect -687 361 -669 395
rect -739 314 -669 361
rect -611 395 -541 411
rect -611 361 -593 395
rect -559 361 -541 395
rect -611 314 -541 361
rect -483 395 -413 411
rect -483 361 -465 395
rect -431 361 -413 395
rect -483 314 -413 361
rect -355 395 -285 411
rect -355 361 -337 395
rect -303 361 -285 395
rect -355 314 -285 361
rect -227 395 -157 411
rect -227 361 -209 395
rect -175 361 -157 395
rect -227 314 -157 361
rect -99 395 -29 411
rect -99 361 -81 395
rect -47 361 -29 395
rect -99 314 -29 361
rect 29 395 99 411
rect 29 361 47 395
rect 81 361 99 395
rect 29 314 99 361
rect 157 395 227 411
rect 157 361 175 395
rect 209 361 227 395
rect 157 314 227 361
rect 285 395 355 411
rect 285 361 303 395
rect 337 361 355 395
rect 285 314 355 361
rect 413 395 483 411
rect 413 361 431 395
rect 465 361 483 395
rect 413 314 483 361
rect 541 395 611 411
rect 541 361 559 395
rect 593 361 611 395
rect 541 314 611 361
rect 669 395 739 411
rect 669 361 687 395
rect 721 361 739 395
rect 669 314 739 361
rect 797 395 867 411
rect 797 361 815 395
rect 849 361 867 395
rect 797 314 867 361
rect 925 395 995 411
rect 925 361 943 395
rect 977 361 995 395
rect 925 314 995 361
rect 1053 395 1123 411
rect 1053 361 1071 395
rect 1105 361 1123 395
rect 1053 314 1123 361
rect 1181 395 1251 411
rect 1181 361 1199 395
rect 1233 361 1251 395
rect 1181 314 1251 361
rect 1309 395 1379 411
rect 1309 361 1327 395
rect 1361 361 1379 395
rect 1309 314 1379 361
rect 1437 395 1507 411
rect 1437 361 1455 395
rect 1489 361 1507 395
rect 1437 314 1507 361
rect 1565 395 1635 411
rect 1565 361 1583 395
rect 1617 361 1635 395
rect 1565 314 1635 361
rect 1693 395 1763 411
rect 1693 361 1711 395
rect 1745 361 1763 395
rect 1693 314 1763 361
rect 1821 395 1891 411
rect 1821 361 1839 395
rect 1873 361 1891 395
rect 1821 314 1891 361
rect 1949 395 2019 411
rect 1949 361 1967 395
rect 2001 361 2019 395
rect 1949 314 2019 361
rect 2077 395 2147 411
rect 2077 361 2095 395
rect 2129 361 2147 395
rect 2077 314 2147 361
rect 2205 395 2275 411
rect 2205 361 2223 395
rect 2257 361 2275 395
rect 2205 314 2275 361
rect 2333 395 2403 411
rect 2333 361 2351 395
rect 2385 361 2403 395
rect 2333 314 2403 361
rect 2461 395 2531 411
rect 2461 361 2479 395
rect 2513 361 2531 395
rect 2461 314 2531 361
rect -2531 -412 -2461 -386
rect -2403 -412 -2333 -386
rect -2275 -412 -2205 -386
rect -2147 -412 -2077 -386
rect -2019 -412 -1949 -386
rect -1891 -412 -1821 -386
rect -1763 -412 -1693 -386
rect -1635 -412 -1565 -386
rect -1507 -412 -1437 -386
rect -1379 -412 -1309 -386
rect -1251 -412 -1181 -386
rect -1123 -412 -1053 -386
rect -995 -412 -925 -386
rect -867 -412 -797 -386
rect -739 -412 -669 -386
rect -611 -412 -541 -386
rect -483 -412 -413 -386
rect -355 -412 -285 -386
rect -227 -412 -157 -386
rect -99 -412 -29 -386
rect 29 -412 99 -386
rect 157 -412 227 -386
rect 285 -412 355 -386
rect 413 -412 483 -386
rect 541 -412 611 -386
rect 669 -412 739 -386
rect 797 -412 867 -386
rect 925 -412 995 -386
rect 1053 -412 1123 -386
rect 1181 -412 1251 -386
rect 1309 -412 1379 -386
rect 1437 -412 1507 -386
rect 1565 -412 1635 -386
rect 1693 -412 1763 -386
rect 1821 -412 1891 -386
rect 1949 -412 2019 -386
rect 2077 -412 2147 -386
rect 2205 -412 2275 -386
rect 2333 -412 2403 -386
rect 2461 -412 2531 -386
<< polycont >>
rect -2513 361 -2479 395
rect -2385 361 -2351 395
rect -2257 361 -2223 395
rect -2129 361 -2095 395
rect -2001 361 -1967 395
rect -1873 361 -1839 395
rect -1745 361 -1711 395
rect -1617 361 -1583 395
rect -1489 361 -1455 395
rect -1361 361 -1327 395
rect -1233 361 -1199 395
rect -1105 361 -1071 395
rect -977 361 -943 395
rect -849 361 -815 395
rect -721 361 -687 395
rect -593 361 -559 395
rect -465 361 -431 395
rect -337 361 -303 395
rect -209 361 -175 395
rect -81 361 -47 395
rect 47 361 81 395
rect 175 361 209 395
rect 303 361 337 395
rect 431 361 465 395
rect 559 361 593 395
rect 687 361 721 395
rect 815 361 849 395
rect 943 361 977 395
rect 1071 361 1105 395
rect 1199 361 1233 395
rect 1327 361 1361 395
rect 1455 361 1489 395
rect 1583 361 1617 395
rect 1711 361 1745 395
rect 1839 361 1873 395
rect 1967 361 2001 395
rect 2095 361 2129 395
rect 2223 361 2257 395
rect 2351 361 2385 395
rect 2479 361 2513 395
<< locali >>
rect -2691 464 -2567 498
rect -2533 464 -2499 498
rect -2465 464 -2431 498
rect -2397 464 -2363 498
rect -2329 464 -2295 498
rect -2261 464 -2227 498
rect -2193 464 -2159 498
rect -2125 464 -2091 498
rect -2057 464 -2023 498
rect -1989 464 -1955 498
rect -1921 464 -1887 498
rect -1853 464 -1819 498
rect -1785 464 -1751 498
rect -1717 464 -1683 498
rect -1649 464 -1615 498
rect -1581 464 -1547 498
rect -1513 464 -1479 498
rect -1445 464 -1411 498
rect -1377 464 -1343 498
rect -1309 464 -1275 498
rect -1241 464 -1207 498
rect -1173 464 -1139 498
rect -1105 464 -1071 498
rect -1037 464 -1003 498
rect -969 464 -935 498
rect -901 464 -867 498
rect -833 464 -799 498
rect -765 464 -731 498
rect -697 464 -663 498
rect -629 464 -595 498
rect -561 464 -527 498
rect -493 464 -459 498
rect -425 464 -391 498
rect -357 464 -323 498
rect -289 464 -255 498
rect -221 464 -187 498
rect -153 464 -119 498
rect -85 464 -51 498
rect -17 464 17 498
rect 51 464 85 498
rect 119 464 153 498
rect 187 464 221 498
rect 255 464 289 498
rect 323 464 357 498
rect 391 464 425 498
rect 459 464 493 498
rect 527 464 561 498
rect 595 464 629 498
rect 663 464 697 498
rect 731 464 765 498
rect 799 464 833 498
rect 867 464 901 498
rect 935 464 969 498
rect 1003 464 1037 498
rect 1071 464 1105 498
rect 1139 464 1173 498
rect 1207 464 1241 498
rect 1275 464 1309 498
rect 1343 464 1377 498
rect 1411 464 1445 498
rect 1479 464 1513 498
rect 1547 464 1581 498
rect 1615 464 1649 498
rect 1683 464 1717 498
rect 1751 464 1785 498
rect 1819 464 1853 498
rect 1887 464 1921 498
rect 1955 464 1989 498
rect 2023 464 2057 498
rect 2091 464 2125 498
rect 2159 464 2193 498
rect 2227 464 2261 498
rect 2295 464 2329 498
rect 2363 464 2397 498
rect 2431 464 2465 498
rect 2499 464 2533 498
rect 2567 464 2691 498
rect -2691 391 -2657 464
rect -2531 361 -2513 395
rect -2479 361 -2461 395
rect -2403 361 -2385 395
rect -2351 361 -2333 395
rect -2275 361 -2257 395
rect -2223 361 -2205 395
rect -2147 361 -2129 395
rect -2095 361 -2077 395
rect -2019 361 -2001 395
rect -1967 361 -1949 395
rect -1891 361 -1873 395
rect -1839 361 -1821 395
rect -1763 361 -1745 395
rect -1711 361 -1693 395
rect -1635 361 -1617 395
rect -1583 361 -1565 395
rect -1507 361 -1489 395
rect -1455 361 -1437 395
rect -1379 361 -1361 395
rect -1327 361 -1309 395
rect -1251 361 -1233 395
rect -1199 361 -1181 395
rect -1123 361 -1105 395
rect -1071 361 -1053 395
rect -995 361 -977 395
rect -943 361 -925 395
rect -867 361 -849 395
rect -815 361 -797 395
rect -739 361 -721 395
rect -687 361 -669 395
rect -611 361 -593 395
rect -559 361 -541 395
rect -483 361 -465 395
rect -431 361 -413 395
rect -355 361 -337 395
rect -303 361 -285 395
rect -227 361 -209 395
rect -175 361 -157 395
rect -99 361 -81 395
rect -47 361 -29 395
rect 29 361 47 395
rect 81 361 99 395
rect 157 361 175 395
rect 209 361 227 395
rect 285 361 303 395
rect 337 361 355 395
rect 413 361 431 395
rect 465 361 483 395
rect 541 361 559 395
rect 593 361 611 395
rect 669 361 687 395
rect 721 361 739 395
rect 797 361 815 395
rect 849 361 867 395
rect 925 361 943 395
rect 977 361 995 395
rect 1053 361 1071 395
rect 1105 361 1123 395
rect 1181 361 1199 395
rect 1233 361 1251 395
rect 1309 361 1327 395
rect 1361 361 1379 395
rect 1437 361 1455 395
rect 1489 361 1507 395
rect 1565 361 1583 395
rect 1617 361 1635 395
rect 1693 361 1711 395
rect 1745 361 1763 395
rect 1821 361 1839 395
rect 1873 361 1891 395
rect 1949 361 1967 395
rect 2001 361 2019 395
rect 2077 361 2095 395
rect 2129 361 2147 395
rect 2205 361 2223 395
rect 2257 361 2275 395
rect 2333 361 2351 395
rect 2385 361 2403 395
rect 2461 361 2479 395
rect 2513 361 2531 395
rect 2657 391 2691 464
rect -2691 323 -2657 357
rect 2657 323 2691 357
rect -2691 255 -2657 289
rect -2691 187 -2657 221
rect -2691 119 -2657 153
rect -2691 51 -2657 85
rect -2691 -17 -2657 17
rect -2691 -85 -2657 -51
rect -2691 -153 -2657 -119
rect -2691 -221 -2657 -187
rect -2691 -289 -2657 -255
rect -2691 -357 -2657 -323
rect -2577 287 -2543 318
rect -2577 219 -2543 235
rect -2577 151 -2543 163
rect -2577 83 -2543 91
rect -2577 15 -2543 19
rect -2577 -91 -2543 -87
rect -2577 -163 -2543 -155
rect -2577 -235 -2543 -223
rect -2577 -307 -2543 -291
rect -2577 -390 -2543 -359
rect -2449 287 -2415 318
rect -2449 219 -2415 235
rect -2449 151 -2415 163
rect -2449 83 -2415 91
rect -2449 15 -2415 19
rect -2449 -91 -2415 -87
rect -2449 -163 -2415 -155
rect -2449 -235 -2415 -223
rect -2449 -307 -2415 -291
rect -2449 -390 -2415 -359
rect -2321 287 -2287 318
rect -2321 219 -2287 235
rect -2321 151 -2287 163
rect -2321 83 -2287 91
rect -2321 15 -2287 19
rect -2321 -91 -2287 -87
rect -2321 -163 -2287 -155
rect -2321 -235 -2287 -223
rect -2321 -307 -2287 -291
rect -2321 -390 -2287 -359
rect -2193 287 -2159 318
rect -2193 219 -2159 235
rect -2193 151 -2159 163
rect -2193 83 -2159 91
rect -2193 15 -2159 19
rect -2193 -91 -2159 -87
rect -2193 -163 -2159 -155
rect -2193 -235 -2159 -223
rect -2193 -307 -2159 -291
rect -2193 -390 -2159 -359
rect -2065 287 -2031 318
rect -2065 219 -2031 235
rect -2065 151 -2031 163
rect -2065 83 -2031 91
rect -2065 15 -2031 19
rect -2065 -91 -2031 -87
rect -2065 -163 -2031 -155
rect -2065 -235 -2031 -223
rect -2065 -307 -2031 -291
rect -2065 -390 -2031 -359
rect -1937 287 -1903 318
rect -1937 219 -1903 235
rect -1937 151 -1903 163
rect -1937 83 -1903 91
rect -1937 15 -1903 19
rect -1937 -91 -1903 -87
rect -1937 -163 -1903 -155
rect -1937 -235 -1903 -223
rect -1937 -307 -1903 -291
rect -1937 -390 -1903 -359
rect -1809 287 -1775 318
rect -1809 219 -1775 235
rect -1809 151 -1775 163
rect -1809 83 -1775 91
rect -1809 15 -1775 19
rect -1809 -91 -1775 -87
rect -1809 -163 -1775 -155
rect -1809 -235 -1775 -223
rect -1809 -307 -1775 -291
rect -1809 -390 -1775 -359
rect -1681 287 -1647 318
rect -1681 219 -1647 235
rect -1681 151 -1647 163
rect -1681 83 -1647 91
rect -1681 15 -1647 19
rect -1681 -91 -1647 -87
rect -1681 -163 -1647 -155
rect -1681 -235 -1647 -223
rect -1681 -307 -1647 -291
rect -1681 -390 -1647 -359
rect -1553 287 -1519 318
rect -1553 219 -1519 235
rect -1553 151 -1519 163
rect -1553 83 -1519 91
rect -1553 15 -1519 19
rect -1553 -91 -1519 -87
rect -1553 -163 -1519 -155
rect -1553 -235 -1519 -223
rect -1553 -307 -1519 -291
rect -1553 -390 -1519 -359
rect -1425 287 -1391 318
rect -1425 219 -1391 235
rect -1425 151 -1391 163
rect -1425 83 -1391 91
rect -1425 15 -1391 19
rect -1425 -91 -1391 -87
rect -1425 -163 -1391 -155
rect -1425 -235 -1391 -223
rect -1425 -307 -1391 -291
rect -1425 -390 -1391 -359
rect -1297 287 -1263 318
rect -1297 219 -1263 235
rect -1297 151 -1263 163
rect -1297 83 -1263 91
rect -1297 15 -1263 19
rect -1297 -91 -1263 -87
rect -1297 -163 -1263 -155
rect -1297 -235 -1263 -223
rect -1297 -307 -1263 -291
rect -1297 -390 -1263 -359
rect -1169 287 -1135 318
rect -1169 219 -1135 235
rect -1169 151 -1135 163
rect -1169 83 -1135 91
rect -1169 15 -1135 19
rect -1169 -91 -1135 -87
rect -1169 -163 -1135 -155
rect -1169 -235 -1135 -223
rect -1169 -307 -1135 -291
rect -1169 -390 -1135 -359
rect -1041 287 -1007 318
rect -1041 219 -1007 235
rect -1041 151 -1007 163
rect -1041 83 -1007 91
rect -1041 15 -1007 19
rect -1041 -91 -1007 -87
rect -1041 -163 -1007 -155
rect -1041 -235 -1007 -223
rect -1041 -307 -1007 -291
rect -1041 -390 -1007 -359
rect -913 287 -879 318
rect -913 219 -879 235
rect -913 151 -879 163
rect -913 83 -879 91
rect -913 15 -879 19
rect -913 -91 -879 -87
rect -913 -163 -879 -155
rect -913 -235 -879 -223
rect -913 -307 -879 -291
rect -913 -390 -879 -359
rect -785 287 -751 318
rect -785 219 -751 235
rect -785 151 -751 163
rect -785 83 -751 91
rect -785 15 -751 19
rect -785 -91 -751 -87
rect -785 -163 -751 -155
rect -785 -235 -751 -223
rect -785 -307 -751 -291
rect -785 -390 -751 -359
rect -657 287 -623 318
rect -657 219 -623 235
rect -657 151 -623 163
rect -657 83 -623 91
rect -657 15 -623 19
rect -657 -91 -623 -87
rect -657 -163 -623 -155
rect -657 -235 -623 -223
rect -657 -307 -623 -291
rect -657 -390 -623 -359
rect -529 287 -495 318
rect -529 219 -495 235
rect -529 151 -495 163
rect -529 83 -495 91
rect -529 15 -495 19
rect -529 -91 -495 -87
rect -529 -163 -495 -155
rect -529 -235 -495 -223
rect -529 -307 -495 -291
rect -529 -390 -495 -359
rect -401 287 -367 318
rect -401 219 -367 235
rect -401 151 -367 163
rect -401 83 -367 91
rect -401 15 -367 19
rect -401 -91 -367 -87
rect -401 -163 -367 -155
rect -401 -235 -367 -223
rect -401 -307 -367 -291
rect -401 -390 -367 -359
rect -273 287 -239 318
rect -273 219 -239 235
rect -273 151 -239 163
rect -273 83 -239 91
rect -273 15 -239 19
rect -273 -91 -239 -87
rect -273 -163 -239 -155
rect -273 -235 -239 -223
rect -273 -307 -239 -291
rect -273 -390 -239 -359
rect -145 287 -111 318
rect -145 219 -111 235
rect -145 151 -111 163
rect -145 83 -111 91
rect -145 15 -111 19
rect -145 -91 -111 -87
rect -145 -163 -111 -155
rect -145 -235 -111 -223
rect -145 -307 -111 -291
rect -145 -390 -111 -359
rect -17 287 17 318
rect -17 219 17 235
rect -17 151 17 163
rect -17 83 17 91
rect -17 15 17 19
rect -17 -91 17 -87
rect -17 -163 17 -155
rect -17 -235 17 -223
rect -17 -307 17 -291
rect -17 -390 17 -359
rect 111 287 145 318
rect 111 219 145 235
rect 111 151 145 163
rect 111 83 145 91
rect 111 15 145 19
rect 111 -91 145 -87
rect 111 -163 145 -155
rect 111 -235 145 -223
rect 111 -307 145 -291
rect 111 -390 145 -359
rect 239 287 273 318
rect 239 219 273 235
rect 239 151 273 163
rect 239 83 273 91
rect 239 15 273 19
rect 239 -91 273 -87
rect 239 -163 273 -155
rect 239 -235 273 -223
rect 239 -307 273 -291
rect 239 -390 273 -359
rect 367 287 401 318
rect 367 219 401 235
rect 367 151 401 163
rect 367 83 401 91
rect 367 15 401 19
rect 367 -91 401 -87
rect 367 -163 401 -155
rect 367 -235 401 -223
rect 367 -307 401 -291
rect 367 -390 401 -359
rect 495 287 529 318
rect 495 219 529 235
rect 495 151 529 163
rect 495 83 529 91
rect 495 15 529 19
rect 495 -91 529 -87
rect 495 -163 529 -155
rect 495 -235 529 -223
rect 495 -307 529 -291
rect 495 -390 529 -359
rect 623 287 657 318
rect 623 219 657 235
rect 623 151 657 163
rect 623 83 657 91
rect 623 15 657 19
rect 623 -91 657 -87
rect 623 -163 657 -155
rect 623 -235 657 -223
rect 623 -307 657 -291
rect 623 -390 657 -359
rect 751 287 785 318
rect 751 219 785 235
rect 751 151 785 163
rect 751 83 785 91
rect 751 15 785 19
rect 751 -91 785 -87
rect 751 -163 785 -155
rect 751 -235 785 -223
rect 751 -307 785 -291
rect 751 -390 785 -359
rect 879 287 913 318
rect 879 219 913 235
rect 879 151 913 163
rect 879 83 913 91
rect 879 15 913 19
rect 879 -91 913 -87
rect 879 -163 913 -155
rect 879 -235 913 -223
rect 879 -307 913 -291
rect 879 -390 913 -359
rect 1007 287 1041 318
rect 1007 219 1041 235
rect 1007 151 1041 163
rect 1007 83 1041 91
rect 1007 15 1041 19
rect 1007 -91 1041 -87
rect 1007 -163 1041 -155
rect 1007 -235 1041 -223
rect 1007 -307 1041 -291
rect 1007 -390 1041 -359
rect 1135 287 1169 318
rect 1135 219 1169 235
rect 1135 151 1169 163
rect 1135 83 1169 91
rect 1135 15 1169 19
rect 1135 -91 1169 -87
rect 1135 -163 1169 -155
rect 1135 -235 1169 -223
rect 1135 -307 1169 -291
rect 1135 -390 1169 -359
rect 1263 287 1297 318
rect 1263 219 1297 235
rect 1263 151 1297 163
rect 1263 83 1297 91
rect 1263 15 1297 19
rect 1263 -91 1297 -87
rect 1263 -163 1297 -155
rect 1263 -235 1297 -223
rect 1263 -307 1297 -291
rect 1263 -390 1297 -359
rect 1391 287 1425 318
rect 1391 219 1425 235
rect 1391 151 1425 163
rect 1391 83 1425 91
rect 1391 15 1425 19
rect 1391 -91 1425 -87
rect 1391 -163 1425 -155
rect 1391 -235 1425 -223
rect 1391 -307 1425 -291
rect 1391 -390 1425 -359
rect 1519 287 1553 318
rect 1519 219 1553 235
rect 1519 151 1553 163
rect 1519 83 1553 91
rect 1519 15 1553 19
rect 1519 -91 1553 -87
rect 1519 -163 1553 -155
rect 1519 -235 1553 -223
rect 1519 -307 1553 -291
rect 1519 -390 1553 -359
rect 1647 287 1681 318
rect 1647 219 1681 235
rect 1647 151 1681 163
rect 1647 83 1681 91
rect 1647 15 1681 19
rect 1647 -91 1681 -87
rect 1647 -163 1681 -155
rect 1647 -235 1681 -223
rect 1647 -307 1681 -291
rect 1647 -390 1681 -359
rect 1775 287 1809 318
rect 1775 219 1809 235
rect 1775 151 1809 163
rect 1775 83 1809 91
rect 1775 15 1809 19
rect 1775 -91 1809 -87
rect 1775 -163 1809 -155
rect 1775 -235 1809 -223
rect 1775 -307 1809 -291
rect 1775 -390 1809 -359
rect 1903 287 1937 318
rect 1903 219 1937 235
rect 1903 151 1937 163
rect 1903 83 1937 91
rect 1903 15 1937 19
rect 1903 -91 1937 -87
rect 1903 -163 1937 -155
rect 1903 -235 1937 -223
rect 1903 -307 1937 -291
rect 1903 -390 1937 -359
rect 2031 287 2065 318
rect 2031 219 2065 235
rect 2031 151 2065 163
rect 2031 83 2065 91
rect 2031 15 2065 19
rect 2031 -91 2065 -87
rect 2031 -163 2065 -155
rect 2031 -235 2065 -223
rect 2031 -307 2065 -291
rect 2031 -390 2065 -359
rect 2159 287 2193 318
rect 2159 219 2193 235
rect 2159 151 2193 163
rect 2159 83 2193 91
rect 2159 15 2193 19
rect 2159 -91 2193 -87
rect 2159 -163 2193 -155
rect 2159 -235 2193 -223
rect 2159 -307 2193 -291
rect 2159 -390 2193 -359
rect 2287 287 2321 318
rect 2287 219 2321 235
rect 2287 151 2321 163
rect 2287 83 2321 91
rect 2287 15 2321 19
rect 2287 -91 2321 -87
rect 2287 -163 2321 -155
rect 2287 -235 2321 -223
rect 2287 -307 2321 -291
rect 2287 -390 2321 -359
rect 2415 287 2449 318
rect 2415 219 2449 235
rect 2415 151 2449 163
rect 2415 83 2449 91
rect 2415 15 2449 19
rect 2415 -91 2449 -87
rect 2415 -163 2449 -155
rect 2415 -235 2449 -223
rect 2415 -307 2449 -291
rect 2415 -390 2449 -359
rect 2543 287 2577 318
rect 2543 219 2577 235
rect 2543 151 2577 163
rect 2543 83 2577 91
rect 2543 15 2577 19
rect 2543 -91 2577 -87
rect 2543 -163 2577 -155
rect 2543 -235 2577 -223
rect 2543 -307 2577 -291
rect 2543 -390 2577 -359
rect 2657 255 2691 289
rect 2657 187 2691 221
rect 2657 119 2691 153
rect 2657 51 2691 85
rect 2657 -17 2691 17
rect 2657 -85 2691 -51
rect 2657 -153 2691 -119
rect 2657 -221 2691 -187
rect 2657 -289 2691 -255
rect 2657 -357 2691 -323
rect -2691 -464 -2657 -391
rect 2657 -464 2691 -391
rect -2691 -498 -2567 -464
rect -2533 -498 -2499 -464
rect -2465 -498 -2431 -464
rect -2397 -498 -2363 -464
rect -2329 -498 -2295 -464
rect -2261 -498 -2227 -464
rect -2193 -498 -2159 -464
rect -2125 -498 -2091 -464
rect -2057 -498 -2023 -464
rect -1989 -498 -1955 -464
rect -1921 -498 -1887 -464
rect -1853 -498 -1819 -464
rect -1785 -498 -1751 -464
rect -1717 -498 -1683 -464
rect -1649 -498 -1615 -464
rect -1581 -498 -1547 -464
rect -1513 -498 -1479 -464
rect -1445 -498 -1411 -464
rect -1377 -498 -1343 -464
rect -1309 -498 -1275 -464
rect -1241 -498 -1207 -464
rect -1173 -498 -1139 -464
rect -1105 -498 -1071 -464
rect -1037 -498 -1003 -464
rect -969 -498 -935 -464
rect -901 -498 -867 -464
rect -833 -498 -799 -464
rect -765 -498 -731 -464
rect -697 -498 -663 -464
rect -629 -498 -595 -464
rect -561 -498 -527 -464
rect -493 -498 -459 -464
rect -425 -498 -391 -464
rect -357 -498 -323 -464
rect -289 -498 -255 -464
rect -221 -498 -187 -464
rect -153 -498 -119 -464
rect -85 -498 -51 -464
rect -17 -498 17 -464
rect 51 -498 85 -464
rect 119 -498 153 -464
rect 187 -498 221 -464
rect 255 -498 289 -464
rect 323 -498 357 -464
rect 391 -498 425 -464
rect 459 -498 493 -464
rect 527 -498 561 -464
rect 595 -498 629 -464
rect 663 -498 697 -464
rect 731 -498 765 -464
rect 799 -498 833 -464
rect 867 -498 901 -464
rect 935 -498 969 -464
rect 1003 -498 1037 -464
rect 1071 -498 1105 -464
rect 1139 -498 1173 -464
rect 1207 -498 1241 -464
rect 1275 -498 1309 -464
rect 1343 -498 1377 -464
rect 1411 -498 1445 -464
rect 1479 -498 1513 -464
rect 1547 -498 1581 -464
rect 1615 -498 1649 -464
rect 1683 -498 1717 -464
rect 1751 -498 1785 -464
rect 1819 -498 1853 -464
rect 1887 -498 1921 -464
rect 1955 -498 1989 -464
rect 2023 -498 2057 -464
rect 2091 -498 2125 -464
rect 2159 -498 2193 -464
rect 2227 -498 2261 -464
rect 2295 -498 2329 -464
rect 2363 -498 2397 -464
rect 2431 -498 2465 -464
rect 2499 -498 2533 -464
rect 2567 -498 2691 -464
<< viali >>
rect -2513 361 -2479 395
rect -2385 361 -2351 395
rect -2257 361 -2223 395
rect -2129 361 -2095 395
rect -2001 361 -1967 395
rect -1873 361 -1839 395
rect -1745 361 -1711 395
rect -1617 361 -1583 395
rect -1489 361 -1455 395
rect -1361 361 -1327 395
rect -1233 361 -1199 395
rect -1105 361 -1071 395
rect -977 361 -943 395
rect -849 361 -815 395
rect -721 361 -687 395
rect -593 361 -559 395
rect -465 361 -431 395
rect -337 361 -303 395
rect -209 361 -175 395
rect -81 361 -47 395
rect 47 361 81 395
rect 175 361 209 395
rect 303 361 337 395
rect 431 361 465 395
rect 559 361 593 395
rect 687 361 721 395
rect 815 361 849 395
rect 943 361 977 395
rect 1071 361 1105 395
rect 1199 361 1233 395
rect 1327 361 1361 395
rect 1455 361 1489 395
rect 1583 361 1617 395
rect 1711 361 1745 395
rect 1839 361 1873 395
rect 1967 361 2001 395
rect 2095 361 2129 395
rect 2223 361 2257 395
rect 2351 361 2385 395
rect 2479 361 2513 395
rect -2577 253 -2543 269
rect -2577 235 -2543 253
rect -2577 185 -2543 197
rect -2577 163 -2543 185
rect -2577 117 -2543 125
rect -2577 91 -2543 117
rect -2577 49 -2543 53
rect -2577 19 -2543 49
rect -2577 -53 -2543 -19
rect -2577 -121 -2543 -91
rect -2577 -125 -2543 -121
rect -2577 -189 -2543 -163
rect -2577 -197 -2543 -189
rect -2577 -257 -2543 -235
rect -2577 -269 -2543 -257
rect -2577 -325 -2543 -307
rect -2577 -341 -2543 -325
rect -2449 253 -2415 269
rect -2449 235 -2415 253
rect -2449 185 -2415 197
rect -2449 163 -2415 185
rect -2449 117 -2415 125
rect -2449 91 -2415 117
rect -2449 49 -2415 53
rect -2449 19 -2415 49
rect -2449 -53 -2415 -19
rect -2449 -121 -2415 -91
rect -2449 -125 -2415 -121
rect -2449 -189 -2415 -163
rect -2449 -197 -2415 -189
rect -2449 -257 -2415 -235
rect -2449 -269 -2415 -257
rect -2449 -325 -2415 -307
rect -2449 -341 -2415 -325
rect -2321 253 -2287 269
rect -2321 235 -2287 253
rect -2321 185 -2287 197
rect -2321 163 -2287 185
rect -2321 117 -2287 125
rect -2321 91 -2287 117
rect -2321 49 -2287 53
rect -2321 19 -2287 49
rect -2321 -53 -2287 -19
rect -2321 -121 -2287 -91
rect -2321 -125 -2287 -121
rect -2321 -189 -2287 -163
rect -2321 -197 -2287 -189
rect -2321 -257 -2287 -235
rect -2321 -269 -2287 -257
rect -2321 -325 -2287 -307
rect -2321 -341 -2287 -325
rect -2193 253 -2159 269
rect -2193 235 -2159 253
rect -2193 185 -2159 197
rect -2193 163 -2159 185
rect -2193 117 -2159 125
rect -2193 91 -2159 117
rect -2193 49 -2159 53
rect -2193 19 -2159 49
rect -2193 -53 -2159 -19
rect -2193 -121 -2159 -91
rect -2193 -125 -2159 -121
rect -2193 -189 -2159 -163
rect -2193 -197 -2159 -189
rect -2193 -257 -2159 -235
rect -2193 -269 -2159 -257
rect -2193 -325 -2159 -307
rect -2193 -341 -2159 -325
rect -2065 253 -2031 269
rect -2065 235 -2031 253
rect -2065 185 -2031 197
rect -2065 163 -2031 185
rect -2065 117 -2031 125
rect -2065 91 -2031 117
rect -2065 49 -2031 53
rect -2065 19 -2031 49
rect -2065 -53 -2031 -19
rect -2065 -121 -2031 -91
rect -2065 -125 -2031 -121
rect -2065 -189 -2031 -163
rect -2065 -197 -2031 -189
rect -2065 -257 -2031 -235
rect -2065 -269 -2031 -257
rect -2065 -325 -2031 -307
rect -2065 -341 -2031 -325
rect -1937 253 -1903 269
rect -1937 235 -1903 253
rect -1937 185 -1903 197
rect -1937 163 -1903 185
rect -1937 117 -1903 125
rect -1937 91 -1903 117
rect -1937 49 -1903 53
rect -1937 19 -1903 49
rect -1937 -53 -1903 -19
rect -1937 -121 -1903 -91
rect -1937 -125 -1903 -121
rect -1937 -189 -1903 -163
rect -1937 -197 -1903 -189
rect -1937 -257 -1903 -235
rect -1937 -269 -1903 -257
rect -1937 -325 -1903 -307
rect -1937 -341 -1903 -325
rect -1809 253 -1775 269
rect -1809 235 -1775 253
rect -1809 185 -1775 197
rect -1809 163 -1775 185
rect -1809 117 -1775 125
rect -1809 91 -1775 117
rect -1809 49 -1775 53
rect -1809 19 -1775 49
rect -1809 -53 -1775 -19
rect -1809 -121 -1775 -91
rect -1809 -125 -1775 -121
rect -1809 -189 -1775 -163
rect -1809 -197 -1775 -189
rect -1809 -257 -1775 -235
rect -1809 -269 -1775 -257
rect -1809 -325 -1775 -307
rect -1809 -341 -1775 -325
rect -1681 253 -1647 269
rect -1681 235 -1647 253
rect -1681 185 -1647 197
rect -1681 163 -1647 185
rect -1681 117 -1647 125
rect -1681 91 -1647 117
rect -1681 49 -1647 53
rect -1681 19 -1647 49
rect -1681 -53 -1647 -19
rect -1681 -121 -1647 -91
rect -1681 -125 -1647 -121
rect -1681 -189 -1647 -163
rect -1681 -197 -1647 -189
rect -1681 -257 -1647 -235
rect -1681 -269 -1647 -257
rect -1681 -325 -1647 -307
rect -1681 -341 -1647 -325
rect -1553 253 -1519 269
rect -1553 235 -1519 253
rect -1553 185 -1519 197
rect -1553 163 -1519 185
rect -1553 117 -1519 125
rect -1553 91 -1519 117
rect -1553 49 -1519 53
rect -1553 19 -1519 49
rect -1553 -53 -1519 -19
rect -1553 -121 -1519 -91
rect -1553 -125 -1519 -121
rect -1553 -189 -1519 -163
rect -1553 -197 -1519 -189
rect -1553 -257 -1519 -235
rect -1553 -269 -1519 -257
rect -1553 -325 -1519 -307
rect -1553 -341 -1519 -325
rect -1425 253 -1391 269
rect -1425 235 -1391 253
rect -1425 185 -1391 197
rect -1425 163 -1391 185
rect -1425 117 -1391 125
rect -1425 91 -1391 117
rect -1425 49 -1391 53
rect -1425 19 -1391 49
rect -1425 -53 -1391 -19
rect -1425 -121 -1391 -91
rect -1425 -125 -1391 -121
rect -1425 -189 -1391 -163
rect -1425 -197 -1391 -189
rect -1425 -257 -1391 -235
rect -1425 -269 -1391 -257
rect -1425 -325 -1391 -307
rect -1425 -341 -1391 -325
rect -1297 253 -1263 269
rect -1297 235 -1263 253
rect -1297 185 -1263 197
rect -1297 163 -1263 185
rect -1297 117 -1263 125
rect -1297 91 -1263 117
rect -1297 49 -1263 53
rect -1297 19 -1263 49
rect -1297 -53 -1263 -19
rect -1297 -121 -1263 -91
rect -1297 -125 -1263 -121
rect -1297 -189 -1263 -163
rect -1297 -197 -1263 -189
rect -1297 -257 -1263 -235
rect -1297 -269 -1263 -257
rect -1297 -325 -1263 -307
rect -1297 -341 -1263 -325
rect -1169 253 -1135 269
rect -1169 235 -1135 253
rect -1169 185 -1135 197
rect -1169 163 -1135 185
rect -1169 117 -1135 125
rect -1169 91 -1135 117
rect -1169 49 -1135 53
rect -1169 19 -1135 49
rect -1169 -53 -1135 -19
rect -1169 -121 -1135 -91
rect -1169 -125 -1135 -121
rect -1169 -189 -1135 -163
rect -1169 -197 -1135 -189
rect -1169 -257 -1135 -235
rect -1169 -269 -1135 -257
rect -1169 -325 -1135 -307
rect -1169 -341 -1135 -325
rect -1041 253 -1007 269
rect -1041 235 -1007 253
rect -1041 185 -1007 197
rect -1041 163 -1007 185
rect -1041 117 -1007 125
rect -1041 91 -1007 117
rect -1041 49 -1007 53
rect -1041 19 -1007 49
rect -1041 -53 -1007 -19
rect -1041 -121 -1007 -91
rect -1041 -125 -1007 -121
rect -1041 -189 -1007 -163
rect -1041 -197 -1007 -189
rect -1041 -257 -1007 -235
rect -1041 -269 -1007 -257
rect -1041 -325 -1007 -307
rect -1041 -341 -1007 -325
rect -913 253 -879 269
rect -913 235 -879 253
rect -913 185 -879 197
rect -913 163 -879 185
rect -913 117 -879 125
rect -913 91 -879 117
rect -913 49 -879 53
rect -913 19 -879 49
rect -913 -53 -879 -19
rect -913 -121 -879 -91
rect -913 -125 -879 -121
rect -913 -189 -879 -163
rect -913 -197 -879 -189
rect -913 -257 -879 -235
rect -913 -269 -879 -257
rect -913 -325 -879 -307
rect -913 -341 -879 -325
rect -785 253 -751 269
rect -785 235 -751 253
rect -785 185 -751 197
rect -785 163 -751 185
rect -785 117 -751 125
rect -785 91 -751 117
rect -785 49 -751 53
rect -785 19 -751 49
rect -785 -53 -751 -19
rect -785 -121 -751 -91
rect -785 -125 -751 -121
rect -785 -189 -751 -163
rect -785 -197 -751 -189
rect -785 -257 -751 -235
rect -785 -269 -751 -257
rect -785 -325 -751 -307
rect -785 -341 -751 -325
rect -657 253 -623 269
rect -657 235 -623 253
rect -657 185 -623 197
rect -657 163 -623 185
rect -657 117 -623 125
rect -657 91 -623 117
rect -657 49 -623 53
rect -657 19 -623 49
rect -657 -53 -623 -19
rect -657 -121 -623 -91
rect -657 -125 -623 -121
rect -657 -189 -623 -163
rect -657 -197 -623 -189
rect -657 -257 -623 -235
rect -657 -269 -623 -257
rect -657 -325 -623 -307
rect -657 -341 -623 -325
rect -529 253 -495 269
rect -529 235 -495 253
rect -529 185 -495 197
rect -529 163 -495 185
rect -529 117 -495 125
rect -529 91 -495 117
rect -529 49 -495 53
rect -529 19 -495 49
rect -529 -53 -495 -19
rect -529 -121 -495 -91
rect -529 -125 -495 -121
rect -529 -189 -495 -163
rect -529 -197 -495 -189
rect -529 -257 -495 -235
rect -529 -269 -495 -257
rect -529 -325 -495 -307
rect -529 -341 -495 -325
rect -401 253 -367 269
rect -401 235 -367 253
rect -401 185 -367 197
rect -401 163 -367 185
rect -401 117 -367 125
rect -401 91 -367 117
rect -401 49 -367 53
rect -401 19 -367 49
rect -401 -53 -367 -19
rect -401 -121 -367 -91
rect -401 -125 -367 -121
rect -401 -189 -367 -163
rect -401 -197 -367 -189
rect -401 -257 -367 -235
rect -401 -269 -367 -257
rect -401 -325 -367 -307
rect -401 -341 -367 -325
rect -273 253 -239 269
rect -273 235 -239 253
rect -273 185 -239 197
rect -273 163 -239 185
rect -273 117 -239 125
rect -273 91 -239 117
rect -273 49 -239 53
rect -273 19 -239 49
rect -273 -53 -239 -19
rect -273 -121 -239 -91
rect -273 -125 -239 -121
rect -273 -189 -239 -163
rect -273 -197 -239 -189
rect -273 -257 -239 -235
rect -273 -269 -239 -257
rect -273 -325 -239 -307
rect -273 -341 -239 -325
rect -145 253 -111 269
rect -145 235 -111 253
rect -145 185 -111 197
rect -145 163 -111 185
rect -145 117 -111 125
rect -145 91 -111 117
rect -145 49 -111 53
rect -145 19 -111 49
rect -145 -53 -111 -19
rect -145 -121 -111 -91
rect -145 -125 -111 -121
rect -145 -189 -111 -163
rect -145 -197 -111 -189
rect -145 -257 -111 -235
rect -145 -269 -111 -257
rect -145 -325 -111 -307
rect -145 -341 -111 -325
rect -17 253 17 269
rect -17 235 17 253
rect -17 185 17 197
rect -17 163 17 185
rect -17 117 17 125
rect -17 91 17 117
rect -17 49 17 53
rect -17 19 17 49
rect -17 -53 17 -19
rect -17 -121 17 -91
rect -17 -125 17 -121
rect -17 -189 17 -163
rect -17 -197 17 -189
rect -17 -257 17 -235
rect -17 -269 17 -257
rect -17 -325 17 -307
rect -17 -341 17 -325
rect 111 253 145 269
rect 111 235 145 253
rect 111 185 145 197
rect 111 163 145 185
rect 111 117 145 125
rect 111 91 145 117
rect 111 49 145 53
rect 111 19 145 49
rect 111 -53 145 -19
rect 111 -121 145 -91
rect 111 -125 145 -121
rect 111 -189 145 -163
rect 111 -197 145 -189
rect 111 -257 145 -235
rect 111 -269 145 -257
rect 111 -325 145 -307
rect 111 -341 145 -325
rect 239 253 273 269
rect 239 235 273 253
rect 239 185 273 197
rect 239 163 273 185
rect 239 117 273 125
rect 239 91 273 117
rect 239 49 273 53
rect 239 19 273 49
rect 239 -53 273 -19
rect 239 -121 273 -91
rect 239 -125 273 -121
rect 239 -189 273 -163
rect 239 -197 273 -189
rect 239 -257 273 -235
rect 239 -269 273 -257
rect 239 -325 273 -307
rect 239 -341 273 -325
rect 367 253 401 269
rect 367 235 401 253
rect 367 185 401 197
rect 367 163 401 185
rect 367 117 401 125
rect 367 91 401 117
rect 367 49 401 53
rect 367 19 401 49
rect 367 -53 401 -19
rect 367 -121 401 -91
rect 367 -125 401 -121
rect 367 -189 401 -163
rect 367 -197 401 -189
rect 367 -257 401 -235
rect 367 -269 401 -257
rect 367 -325 401 -307
rect 367 -341 401 -325
rect 495 253 529 269
rect 495 235 529 253
rect 495 185 529 197
rect 495 163 529 185
rect 495 117 529 125
rect 495 91 529 117
rect 495 49 529 53
rect 495 19 529 49
rect 495 -53 529 -19
rect 495 -121 529 -91
rect 495 -125 529 -121
rect 495 -189 529 -163
rect 495 -197 529 -189
rect 495 -257 529 -235
rect 495 -269 529 -257
rect 495 -325 529 -307
rect 495 -341 529 -325
rect 623 253 657 269
rect 623 235 657 253
rect 623 185 657 197
rect 623 163 657 185
rect 623 117 657 125
rect 623 91 657 117
rect 623 49 657 53
rect 623 19 657 49
rect 623 -53 657 -19
rect 623 -121 657 -91
rect 623 -125 657 -121
rect 623 -189 657 -163
rect 623 -197 657 -189
rect 623 -257 657 -235
rect 623 -269 657 -257
rect 623 -325 657 -307
rect 623 -341 657 -325
rect 751 253 785 269
rect 751 235 785 253
rect 751 185 785 197
rect 751 163 785 185
rect 751 117 785 125
rect 751 91 785 117
rect 751 49 785 53
rect 751 19 785 49
rect 751 -53 785 -19
rect 751 -121 785 -91
rect 751 -125 785 -121
rect 751 -189 785 -163
rect 751 -197 785 -189
rect 751 -257 785 -235
rect 751 -269 785 -257
rect 751 -325 785 -307
rect 751 -341 785 -325
rect 879 253 913 269
rect 879 235 913 253
rect 879 185 913 197
rect 879 163 913 185
rect 879 117 913 125
rect 879 91 913 117
rect 879 49 913 53
rect 879 19 913 49
rect 879 -53 913 -19
rect 879 -121 913 -91
rect 879 -125 913 -121
rect 879 -189 913 -163
rect 879 -197 913 -189
rect 879 -257 913 -235
rect 879 -269 913 -257
rect 879 -325 913 -307
rect 879 -341 913 -325
rect 1007 253 1041 269
rect 1007 235 1041 253
rect 1007 185 1041 197
rect 1007 163 1041 185
rect 1007 117 1041 125
rect 1007 91 1041 117
rect 1007 49 1041 53
rect 1007 19 1041 49
rect 1007 -53 1041 -19
rect 1007 -121 1041 -91
rect 1007 -125 1041 -121
rect 1007 -189 1041 -163
rect 1007 -197 1041 -189
rect 1007 -257 1041 -235
rect 1007 -269 1041 -257
rect 1007 -325 1041 -307
rect 1007 -341 1041 -325
rect 1135 253 1169 269
rect 1135 235 1169 253
rect 1135 185 1169 197
rect 1135 163 1169 185
rect 1135 117 1169 125
rect 1135 91 1169 117
rect 1135 49 1169 53
rect 1135 19 1169 49
rect 1135 -53 1169 -19
rect 1135 -121 1169 -91
rect 1135 -125 1169 -121
rect 1135 -189 1169 -163
rect 1135 -197 1169 -189
rect 1135 -257 1169 -235
rect 1135 -269 1169 -257
rect 1135 -325 1169 -307
rect 1135 -341 1169 -325
rect 1263 253 1297 269
rect 1263 235 1297 253
rect 1263 185 1297 197
rect 1263 163 1297 185
rect 1263 117 1297 125
rect 1263 91 1297 117
rect 1263 49 1297 53
rect 1263 19 1297 49
rect 1263 -53 1297 -19
rect 1263 -121 1297 -91
rect 1263 -125 1297 -121
rect 1263 -189 1297 -163
rect 1263 -197 1297 -189
rect 1263 -257 1297 -235
rect 1263 -269 1297 -257
rect 1263 -325 1297 -307
rect 1263 -341 1297 -325
rect 1391 253 1425 269
rect 1391 235 1425 253
rect 1391 185 1425 197
rect 1391 163 1425 185
rect 1391 117 1425 125
rect 1391 91 1425 117
rect 1391 49 1425 53
rect 1391 19 1425 49
rect 1391 -53 1425 -19
rect 1391 -121 1425 -91
rect 1391 -125 1425 -121
rect 1391 -189 1425 -163
rect 1391 -197 1425 -189
rect 1391 -257 1425 -235
rect 1391 -269 1425 -257
rect 1391 -325 1425 -307
rect 1391 -341 1425 -325
rect 1519 253 1553 269
rect 1519 235 1553 253
rect 1519 185 1553 197
rect 1519 163 1553 185
rect 1519 117 1553 125
rect 1519 91 1553 117
rect 1519 49 1553 53
rect 1519 19 1553 49
rect 1519 -53 1553 -19
rect 1519 -121 1553 -91
rect 1519 -125 1553 -121
rect 1519 -189 1553 -163
rect 1519 -197 1553 -189
rect 1519 -257 1553 -235
rect 1519 -269 1553 -257
rect 1519 -325 1553 -307
rect 1519 -341 1553 -325
rect 1647 253 1681 269
rect 1647 235 1681 253
rect 1647 185 1681 197
rect 1647 163 1681 185
rect 1647 117 1681 125
rect 1647 91 1681 117
rect 1647 49 1681 53
rect 1647 19 1681 49
rect 1647 -53 1681 -19
rect 1647 -121 1681 -91
rect 1647 -125 1681 -121
rect 1647 -189 1681 -163
rect 1647 -197 1681 -189
rect 1647 -257 1681 -235
rect 1647 -269 1681 -257
rect 1647 -325 1681 -307
rect 1647 -341 1681 -325
rect 1775 253 1809 269
rect 1775 235 1809 253
rect 1775 185 1809 197
rect 1775 163 1809 185
rect 1775 117 1809 125
rect 1775 91 1809 117
rect 1775 49 1809 53
rect 1775 19 1809 49
rect 1775 -53 1809 -19
rect 1775 -121 1809 -91
rect 1775 -125 1809 -121
rect 1775 -189 1809 -163
rect 1775 -197 1809 -189
rect 1775 -257 1809 -235
rect 1775 -269 1809 -257
rect 1775 -325 1809 -307
rect 1775 -341 1809 -325
rect 1903 253 1937 269
rect 1903 235 1937 253
rect 1903 185 1937 197
rect 1903 163 1937 185
rect 1903 117 1937 125
rect 1903 91 1937 117
rect 1903 49 1937 53
rect 1903 19 1937 49
rect 1903 -53 1937 -19
rect 1903 -121 1937 -91
rect 1903 -125 1937 -121
rect 1903 -189 1937 -163
rect 1903 -197 1937 -189
rect 1903 -257 1937 -235
rect 1903 -269 1937 -257
rect 1903 -325 1937 -307
rect 1903 -341 1937 -325
rect 2031 253 2065 269
rect 2031 235 2065 253
rect 2031 185 2065 197
rect 2031 163 2065 185
rect 2031 117 2065 125
rect 2031 91 2065 117
rect 2031 49 2065 53
rect 2031 19 2065 49
rect 2031 -53 2065 -19
rect 2031 -121 2065 -91
rect 2031 -125 2065 -121
rect 2031 -189 2065 -163
rect 2031 -197 2065 -189
rect 2031 -257 2065 -235
rect 2031 -269 2065 -257
rect 2031 -325 2065 -307
rect 2031 -341 2065 -325
rect 2159 253 2193 269
rect 2159 235 2193 253
rect 2159 185 2193 197
rect 2159 163 2193 185
rect 2159 117 2193 125
rect 2159 91 2193 117
rect 2159 49 2193 53
rect 2159 19 2193 49
rect 2159 -53 2193 -19
rect 2159 -121 2193 -91
rect 2159 -125 2193 -121
rect 2159 -189 2193 -163
rect 2159 -197 2193 -189
rect 2159 -257 2193 -235
rect 2159 -269 2193 -257
rect 2159 -325 2193 -307
rect 2159 -341 2193 -325
rect 2287 253 2321 269
rect 2287 235 2321 253
rect 2287 185 2321 197
rect 2287 163 2321 185
rect 2287 117 2321 125
rect 2287 91 2321 117
rect 2287 49 2321 53
rect 2287 19 2321 49
rect 2287 -53 2321 -19
rect 2287 -121 2321 -91
rect 2287 -125 2321 -121
rect 2287 -189 2321 -163
rect 2287 -197 2321 -189
rect 2287 -257 2321 -235
rect 2287 -269 2321 -257
rect 2287 -325 2321 -307
rect 2287 -341 2321 -325
rect 2415 253 2449 269
rect 2415 235 2449 253
rect 2415 185 2449 197
rect 2415 163 2449 185
rect 2415 117 2449 125
rect 2415 91 2449 117
rect 2415 49 2449 53
rect 2415 19 2449 49
rect 2415 -53 2449 -19
rect 2415 -121 2449 -91
rect 2415 -125 2449 -121
rect 2415 -189 2449 -163
rect 2415 -197 2449 -189
rect 2415 -257 2449 -235
rect 2415 -269 2449 -257
rect 2415 -325 2449 -307
rect 2415 -341 2449 -325
rect 2543 253 2577 269
rect 2543 235 2577 253
rect 2543 185 2577 197
rect 2543 163 2577 185
rect 2543 117 2577 125
rect 2543 91 2577 117
rect 2543 49 2577 53
rect 2543 19 2577 49
rect 2543 -53 2577 -19
rect 2543 -121 2577 -91
rect 2543 -125 2577 -121
rect 2543 -189 2577 -163
rect 2543 -197 2577 -189
rect 2543 -257 2577 -235
rect 2543 -269 2577 -257
rect 2543 -325 2577 -307
rect 2543 -341 2577 -325
<< metal1 >>
rect -2527 395 -2465 401
rect -2527 361 -2513 395
rect -2479 361 -2465 395
rect -2527 355 -2465 361
rect -2399 395 -2337 401
rect -2399 361 -2385 395
rect -2351 361 -2337 395
rect -2399 355 -2337 361
rect -2271 395 -2209 401
rect -2271 361 -2257 395
rect -2223 361 -2209 395
rect -2271 355 -2209 361
rect -2143 395 -2081 401
rect -2143 361 -2129 395
rect -2095 361 -2081 395
rect -2143 355 -2081 361
rect -2015 395 -1953 401
rect -2015 361 -2001 395
rect -1967 361 -1953 395
rect -2015 355 -1953 361
rect -1887 395 -1825 401
rect -1887 361 -1873 395
rect -1839 361 -1825 395
rect -1887 355 -1825 361
rect -1759 395 -1697 401
rect -1759 361 -1745 395
rect -1711 361 -1697 395
rect -1759 355 -1697 361
rect -1631 395 -1569 401
rect -1631 361 -1617 395
rect -1583 361 -1569 395
rect -1631 355 -1569 361
rect -1503 395 -1441 401
rect -1503 361 -1489 395
rect -1455 361 -1441 395
rect -1503 355 -1441 361
rect -1375 395 -1313 401
rect -1375 361 -1361 395
rect -1327 361 -1313 395
rect -1375 355 -1313 361
rect -1247 395 -1185 401
rect -1247 361 -1233 395
rect -1199 361 -1185 395
rect -1247 355 -1185 361
rect -1119 395 -1057 401
rect -1119 361 -1105 395
rect -1071 361 -1057 395
rect -1119 355 -1057 361
rect -991 395 -929 401
rect -991 361 -977 395
rect -943 361 -929 395
rect -991 355 -929 361
rect -863 395 -801 401
rect -863 361 -849 395
rect -815 361 -801 395
rect -863 355 -801 361
rect -735 395 -673 401
rect -735 361 -721 395
rect -687 361 -673 395
rect -735 355 -673 361
rect -607 395 -545 401
rect -607 361 -593 395
rect -559 361 -545 395
rect -607 355 -545 361
rect -479 395 -417 401
rect -479 361 -465 395
rect -431 361 -417 395
rect -479 355 -417 361
rect -351 395 -289 401
rect -351 361 -337 395
rect -303 361 -289 395
rect -351 355 -289 361
rect -223 395 -161 401
rect -223 361 -209 395
rect -175 361 -161 395
rect -223 355 -161 361
rect -95 395 -33 401
rect -95 361 -81 395
rect -47 361 -33 395
rect -95 355 -33 361
rect 33 395 95 401
rect 33 361 47 395
rect 81 361 95 395
rect 33 355 95 361
rect 161 395 223 401
rect 161 361 175 395
rect 209 361 223 395
rect 161 355 223 361
rect 289 395 351 401
rect 289 361 303 395
rect 337 361 351 395
rect 289 355 351 361
rect 417 395 479 401
rect 417 361 431 395
rect 465 361 479 395
rect 417 355 479 361
rect 545 395 607 401
rect 545 361 559 395
rect 593 361 607 395
rect 545 355 607 361
rect 673 395 735 401
rect 673 361 687 395
rect 721 361 735 395
rect 673 355 735 361
rect 801 395 863 401
rect 801 361 815 395
rect 849 361 863 395
rect 801 355 863 361
rect 929 395 991 401
rect 929 361 943 395
rect 977 361 991 395
rect 929 355 991 361
rect 1057 395 1119 401
rect 1057 361 1071 395
rect 1105 361 1119 395
rect 1057 355 1119 361
rect 1185 395 1247 401
rect 1185 361 1199 395
rect 1233 361 1247 395
rect 1185 355 1247 361
rect 1313 395 1375 401
rect 1313 361 1327 395
rect 1361 361 1375 395
rect 1313 355 1375 361
rect 1441 395 1503 401
rect 1441 361 1455 395
rect 1489 361 1503 395
rect 1441 355 1503 361
rect 1569 395 1631 401
rect 1569 361 1583 395
rect 1617 361 1631 395
rect 1569 355 1631 361
rect 1697 395 1759 401
rect 1697 361 1711 395
rect 1745 361 1759 395
rect 1697 355 1759 361
rect 1825 395 1887 401
rect 1825 361 1839 395
rect 1873 361 1887 395
rect 1825 355 1887 361
rect 1953 395 2015 401
rect 1953 361 1967 395
rect 2001 361 2015 395
rect 1953 355 2015 361
rect 2081 395 2143 401
rect 2081 361 2095 395
rect 2129 361 2143 395
rect 2081 355 2143 361
rect 2209 395 2271 401
rect 2209 361 2223 395
rect 2257 361 2271 395
rect 2209 355 2271 361
rect 2337 395 2399 401
rect 2337 361 2351 395
rect 2385 361 2399 395
rect 2337 355 2399 361
rect 2465 395 2527 401
rect 2465 361 2479 395
rect 2513 361 2527 395
rect 2465 355 2527 361
rect -2583 269 -2537 314
rect -2583 235 -2577 269
rect -2543 235 -2537 269
rect -2583 197 -2537 235
rect -2583 163 -2577 197
rect -2543 163 -2537 197
rect -2583 125 -2537 163
rect -2583 91 -2577 125
rect -2543 91 -2537 125
rect -2583 53 -2537 91
rect -2583 19 -2577 53
rect -2543 19 -2537 53
rect -2583 -19 -2537 19
rect -2583 -53 -2577 -19
rect -2543 -53 -2537 -19
rect -2583 -91 -2537 -53
rect -2583 -125 -2577 -91
rect -2543 -125 -2537 -91
rect -2583 -163 -2537 -125
rect -2583 -197 -2577 -163
rect -2543 -197 -2537 -163
rect -2583 -235 -2537 -197
rect -2583 -269 -2577 -235
rect -2543 -269 -2537 -235
rect -2583 -307 -2537 -269
rect -2583 -341 -2577 -307
rect -2543 -341 -2537 -307
rect -2583 -386 -2537 -341
rect -2455 269 -2409 314
rect -2455 235 -2449 269
rect -2415 235 -2409 269
rect -2455 197 -2409 235
rect -2455 163 -2449 197
rect -2415 163 -2409 197
rect -2455 125 -2409 163
rect -2455 91 -2449 125
rect -2415 91 -2409 125
rect -2455 53 -2409 91
rect -2455 19 -2449 53
rect -2415 19 -2409 53
rect -2455 -19 -2409 19
rect -2455 -53 -2449 -19
rect -2415 -53 -2409 -19
rect -2455 -91 -2409 -53
rect -2455 -125 -2449 -91
rect -2415 -125 -2409 -91
rect -2455 -163 -2409 -125
rect -2455 -197 -2449 -163
rect -2415 -197 -2409 -163
rect -2455 -235 -2409 -197
rect -2455 -269 -2449 -235
rect -2415 -269 -2409 -235
rect -2455 -307 -2409 -269
rect -2455 -341 -2449 -307
rect -2415 -341 -2409 -307
rect -2455 -386 -2409 -341
rect -2327 269 -2281 314
rect -2327 235 -2321 269
rect -2287 235 -2281 269
rect -2327 197 -2281 235
rect -2327 163 -2321 197
rect -2287 163 -2281 197
rect -2327 125 -2281 163
rect -2327 91 -2321 125
rect -2287 91 -2281 125
rect -2327 53 -2281 91
rect -2327 19 -2321 53
rect -2287 19 -2281 53
rect -2327 -19 -2281 19
rect -2327 -53 -2321 -19
rect -2287 -53 -2281 -19
rect -2327 -91 -2281 -53
rect -2327 -125 -2321 -91
rect -2287 -125 -2281 -91
rect -2327 -163 -2281 -125
rect -2327 -197 -2321 -163
rect -2287 -197 -2281 -163
rect -2327 -235 -2281 -197
rect -2327 -269 -2321 -235
rect -2287 -269 -2281 -235
rect -2327 -307 -2281 -269
rect -2327 -341 -2321 -307
rect -2287 -341 -2281 -307
rect -2327 -386 -2281 -341
rect -2199 269 -2153 314
rect -2199 235 -2193 269
rect -2159 235 -2153 269
rect -2199 197 -2153 235
rect -2199 163 -2193 197
rect -2159 163 -2153 197
rect -2199 125 -2153 163
rect -2199 91 -2193 125
rect -2159 91 -2153 125
rect -2199 53 -2153 91
rect -2199 19 -2193 53
rect -2159 19 -2153 53
rect -2199 -19 -2153 19
rect -2199 -53 -2193 -19
rect -2159 -53 -2153 -19
rect -2199 -91 -2153 -53
rect -2199 -125 -2193 -91
rect -2159 -125 -2153 -91
rect -2199 -163 -2153 -125
rect -2199 -197 -2193 -163
rect -2159 -197 -2153 -163
rect -2199 -235 -2153 -197
rect -2199 -269 -2193 -235
rect -2159 -269 -2153 -235
rect -2199 -307 -2153 -269
rect -2199 -341 -2193 -307
rect -2159 -341 -2153 -307
rect -2199 -386 -2153 -341
rect -2071 269 -2025 314
rect -2071 235 -2065 269
rect -2031 235 -2025 269
rect -2071 197 -2025 235
rect -2071 163 -2065 197
rect -2031 163 -2025 197
rect -2071 125 -2025 163
rect -2071 91 -2065 125
rect -2031 91 -2025 125
rect -2071 53 -2025 91
rect -2071 19 -2065 53
rect -2031 19 -2025 53
rect -2071 -19 -2025 19
rect -2071 -53 -2065 -19
rect -2031 -53 -2025 -19
rect -2071 -91 -2025 -53
rect -2071 -125 -2065 -91
rect -2031 -125 -2025 -91
rect -2071 -163 -2025 -125
rect -2071 -197 -2065 -163
rect -2031 -197 -2025 -163
rect -2071 -235 -2025 -197
rect -2071 -269 -2065 -235
rect -2031 -269 -2025 -235
rect -2071 -307 -2025 -269
rect -2071 -341 -2065 -307
rect -2031 -341 -2025 -307
rect -2071 -386 -2025 -341
rect -1943 269 -1897 314
rect -1943 235 -1937 269
rect -1903 235 -1897 269
rect -1943 197 -1897 235
rect -1943 163 -1937 197
rect -1903 163 -1897 197
rect -1943 125 -1897 163
rect -1943 91 -1937 125
rect -1903 91 -1897 125
rect -1943 53 -1897 91
rect -1943 19 -1937 53
rect -1903 19 -1897 53
rect -1943 -19 -1897 19
rect -1943 -53 -1937 -19
rect -1903 -53 -1897 -19
rect -1943 -91 -1897 -53
rect -1943 -125 -1937 -91
rect -1903 -125 -1897 -91
rect -1943 -163 -1897 -125
rect -1943 -197 -1937 -163
rect -1903 -197 -1897 -163
rect -1943 -235 -1897 -197
rect -1943 -269 -1937 -235
rect -1903 -269 -1897 -235
rect -1943 -307 -1897 -269
rect -1943 -341 -1937 -307
rect -1903 -341 -1897 -307
rect -1943 -386 -1897 -341
rect -1815 269 -1769 314
rect -1815 235 -1809 269
rect -1775 235 -1769 269
rect -1815 197 -1769 235
rect -1815 163 -1809 197
rect -1775 163 -1769 197
rect -1815 125 -1769 163
rect -1815 91 -1809 125
rect -1775 91 -1769 125
rect -1815 53 -1769 91
rect -1815 19 -1809 53
rect -1775 19 -1769 53
rect -1815 -19 -1769 19
rect -1815 -53 -1809 -19
rect -1775 -53 -1769 -19
rect -1815 -91 -1769 -53
rect -1815 -125 -1809 -91
rect -1775 -125 -1769 -91
rect -1815 -163 -1769 -125
rect -1815 -197 -1809 -163
rect -1775 -197 -1769 -163
rect -1815 -235 -1769 -197
rect -1815 -269 -1809 -235
rect -1775 -269 -1769 -235
rect -1815 -307 -1769 -269
rect -1815 -341 -1809 -307
rect -1775 -341 -1769 -307
rect -1815 -386 -1769 -341
rect -1687 269 -1641 314
rect -1687 235 -1681 269
rect -1647 235 -1641 269
rect -1687 197 -1641 235
rect -1687 163 -1681 197
rect -1647 163 -1641 197
rect -1687 125 -1641 163
rect -1687 91 -1681 125
rect -1647 91 -1641 125
rect -1687 53 -1641 91
rect -1687 19 -1681 53
rect -1647 19 -1641 53
rect -1687 -19 -1641 19
rect -1687 -53 -1681 -19
rect -1647 -53 -1641 -19
rect -1687 -91 -1641 -53
rect -1687 -125 -1681 -91
rect -1647 -125 -1641 -91
rect -1687 -163 -1641 -125
rect -1687 -197 -1681 -163
rect -1647 -197 -1641 -163
rect -1687 -235 -1641 -197
rect -1687 -269 -1681 -235
rect -1647 -269 -1641 -235
rect -1687 -307 -1641 -269
rect -1687 -341 -1681 -307
rect -1647 -341 -1641 -307
rect -1687 -386 -1641 -341
rect -1559 269 -1513 314
rect -1559 235 -1553 269
rect -1519 235 -1513 269
rect -1559 197 -1513 235
rect -1559 163 -1553 197
rect -1519 163 -1513 197
rect -1559 125 -1513 163
rect -1559 91 -1553 125
rect -1519 91 -1513 125
rect -1559 53 -1513 91
rect -1559 19 -1553 53
rect -1519 19 -1513 53
rect -1559 -19 -1513 19
rect -1559 -53 -1553 -19
rect -1519 -53 -1513 -19
rect -1559 -91 -1513 -53
rect -1559 -125 -1553 -91
rect -1519 -125 -1513 -91
rect -1559 -163 -1513 -125
rect -1559 -197 -1553 -163
rect -1519 -197 -1513 -163
rect -1559 -235 -1513 -197
rect -1559 -269 -1553 -235
rect -1519 -269 -1513 -235
rect -1559 -307 -1513 -269
rect -1559 -341 -1553 -307
rect -1519 -341 -1513 -307
rect -1559 -386 -1513 -341
rect -1431 269 -1385 314
rect -1431 235 -1425 269
rect -1391 235 -1385 269
rect -1431 197 -1385 235
rect -1431 163 -1425 197
rect -1391 163 -1385 197
rect -1431 125 -1385 163
rect -1431 91 -1425 125
rect -1391 91 -1385 125
rect -1431 53 -1385 91
rect -1431 19 -1425 53
rect -1391 19 -1385 53
rect -1431 -19 -1385 19
rect -1431 -53 -1425 -19
rect -1391 -53 -1385 -19
rect -1431 -91 -1385 -53
rect -1431 -125 -1425 -91
rect -1391 -125 -1385 -91
rect -1431 -163 -1385 -125
rect -1431 -197 -1425 -163
rect -1391 -197 -1385 -163
rect -1431 -235 -1385 -197
rect -1431 -269 -1425 -235
rect -1391 -269 -1385 -235
rect -1431 -307 -1385 -269
rect -1431 -341 -1425 -307
rect -1391 -341 -1385 -307
rect -1431 -386 -1385 -341
rect -1303 269 -1257 314
rect -1303 235 -1297 269
rect -1263 235 -1257 269
rect -1303 197 -1257 235
rect -1303 163 -1297 197
rect -1263 163 -1257 197
rect -1303 125 -1257 163
rect -1303 91 -1297 125
rect -1263 91 -1257 125
rect -1303 53 -1257 91
rect -1303 19 -1297 53
rect -1263 19 -1257 53
rect -1303 -19 -1257 19
rect -1303 -53 -1297 -19
rect -1263 -53 -1257 -19
rect -1303 -91 -1257 -53
rect -1303 -125 -1297 -91
rect -1263 -125 -1257 -91
rect -1303 -163 -1257 -125
rect -1303 -197 -1297 -163
rect -1263 -197 -1257 -163
rect -1303 -235 -1257 -197
rect -1303 -269 -1297 -235
rect -1263 -269 -1257 -235
rect -1303 -307 -1257 -269
rect -1303 -341 -1297 -307
rect -1263 -341 -1257 -307
rect -1303 -386 -1257 -341
rect -1175 269 -1129 314
rect -1175 235 -1169 269
rect -1135 235 -1129 269
rect -1175 197 -1129 235
rect -1175 163 -1169 197
rect -1135 163 -1129 197
rect -1175 125 -1129 163
rect -1175 91 -1169 125
rect -1135 91 -1129 125
rect -1175 53 -1129 91
rect -1175 19 -1169 53
rect -1135 19 -1129 53
rect -1175 -19 -1129 19
rect -1175 -53 -1169 -19
rect -1135 -53 -1129 -19
rect -1175 -91 -1129 -53
rect -1175 -125 -1169 -91
rect -1135 -125 -1129 -91
rect -1175 -163 -1129 -125
rect -1175 -197 -1169 -163
rect -1135 -197 -1129 -163
rect -1175 -235 -1129 -197
rect -1175 -269 -1169 -235
rect -1135 -269 -1129 -235
rect -1175 -307 -1129 -269
rect -1175 -341 -1169 -307
rect -1135 -341 -1129 -307
rect -1175 -386 -1129 -341
rect -1047 269 -1001 314
rect -1047 235 -1041 269
rect -1007 235 -1001 269
rect -1047 197 -1001 235
rect -1047 163 -1041 197
rect -1007 163 -1001 197
rect -1047 125 -1001 163
rect -1047 91 -1041 125
rect -1007 91 -1001 125
rect -1047 53 -1001 91
rect -1047 19 -1041 53
rect -1007 19 -1001 53
rect -1047 -19 -1001 19
rect -1047 -53 -1041 -19
rect -1007 -53 -1001 -19
rect -1047 -91 -1001 -53
rect -1047 -125 -1041 -91
rect -1007 -125 -1001 -91
rect -1047 -163 -1001 -125
rect -1047 -197 -1041 -163
rect -1007 -197 -1001 -163
rect -1047 -235 -1001 -197
rect -1047 -269 -1041 -235
rect -1007 -269 -1001 -235
rect -1047 -307 -1001 -269
rect -1047 -341 -1041 -307
rect -1007 -341 -1001 -307
rect -1047 -386 -1001 -341
rect -919 269 -873 314
rect -919 235 -913 269
rect -879 235 -873 269
rect -919 197 -873 235
rect -919 163 -913 197
rect -879 163 -873 197
rect -919 125 -873 163
rect -919 91 -913 125
rect -879 91 -873 125
rect -919 53 -873 91
rect -919 19 -913 53
rect -879 19 -873 53
rect -919 -19 -873 19
rect -919 -53 -913 -19
rect -879 -53 -873 -19
rect -919 -91 -873 -53
rect -919 -125 -913 -91
rect -879 -125 -873 -91
rect -919 -163 -873 -125
rect -919 -197 -913 -163
rect -879 -197 -873 -163
rect -919 -235 -873 -197
rect -919 -269 -913 -235
rect -879 -269 -873 -235
rect -919 -307 -873 -269
rect -919 -341 -913 -307
rect -879 -341 -873 -307
rect -919 -386 -873 -341
rect -791 269 -745 314
rect -791 235 -785 269
rect -751 235 -745 269
rect -791 197 -745 235
rect -791 163 -785 197
rect -751 163 -745 197
rect -791 125 -745 163
rect -791 91 -785 125
rect -751 91 -745 125
rect -791 53 -745 91
rect -791 19 -785 53
rect -751 19 -745 53
rect -791 -19 -745 19
rect -791 -53 -785 -19
rect -751 -53 -745 -19
rect -791 -91 -745 -53
rect -791 -125 -785 -91
rect -751 -125 -745 -91
rect -791 -163 -745 -125
rect -791 -197 -785 -163
rect -751 -197 -745 -163
rect -791 -235 -745 -197
rect -791 -269 -785 -235
rect -751 -269 -745 -235
rect -791 -307 -745 -269
rect -791 -341 -785 -307
rect -751 -341 -745 -307
rect -791 -386 -745 -341
rect -663 269 -617 314
rect -663 235 -657 269
rect -623 235 -617 269
rect -663 197 -617 235
rect -663 163 -657 197
rect -623 163 -617 197
rect -663 125 -617 163
rect -663 91 -657 125
rect -623 91 -617 125
rect -663 53 -617 91
rect -663 19 -657 53
rect -623 19 -617 53
rect -663 -19 -617 19
rect -663 -53 -657 -19
rect -623 -53 -617 -19
rect -663 -91 -617 -53
rect -663 -125 -657 -91
rect -623 -125 -617 -91
rect -663 -163 -617 -125
rect -663 -197 -657 -163
rect -623 -197 -617 -163
rect -663 -235 -617 -197
rect -663 -269 -657 -235
rect -623 -269 -617 -235
rect -663 -307 -617 -269
rect -663 -341 -657 -307
rect -623 -341 -617 -307
rect -663 -386 -617 -341
rect -535 269 -489 314
rect -535 235 -529 269
rect -495 235 -489 269
rect -535 197 -489 235
rect -535 163 -529 197
rect -495 163 -489 197
rect -535 125 -489 163
rect -535 91 -529 125
rect -495 91 -489 125
rect -535 53 -489 91
rect -535 19 -529 53
rect -495 19 -489 53
rect -535 -19 -489 19
rect -535 -53 -529 -19
rect -495 -53 -489 -19
rect -535 -91 -489 -53
rect -535 -125 -529 -91
rect -495 -125 -489 -91
rect -535 -163 -489 -125
rect -535 -197 -529 -163
rect -495 -197 -489 -163
rect -535 -235 -489 -197
rect -535 -269 -529 -235
rect -495 -269 -489 -235
rect -535 -307 -489 -269
rect -535 -341 -529 -307
rect -495 -341 -489 -307
rect -535 -386 -489 -341
rect -407 269 -361 314
rect -407 235 -401 269
rect -367 235 -361 269
rect -407 197 -361 235
rect -407 163 -401 197
rect -367 163 -361 197
rect -407 125 -361 163
rect -407 91 -401 125
rect -367 91 -361 125
rect -407 53 -361 91
rect -407 19 -401 53
rect -367 19 -361 53
rect -407 -19 -361 19
rect -407 -53 -401 -19
rect -367 -53 -361 -19
rect -407 -91 -361 -53
rect -407 -125 -401 -91
rect -367 -125 -361 -91
rect -407 -163 -361 -125
rect -407 -197 -401 -163
rect -367 -197 -361 -163
rect -407 -235 -361 -197
rect -407 -269 -401 -235
rect -367 -269 -361 -235
rect -407 -307 -361 -269
rect -407 -341 -401 -307
rect -367 -341 -361 -307
rect -407 -386 -361 -341
rect -279 269 -233 314
rect -279 235 -273 269
rect -239 235 -233 269
rect -279 197 -233 235
rect -279 163 -273 197
rect -239 163 -233 197
rect -279 125 -233 163
rect -279 91 -273 125
rect -239 91 -233 125
rect -279 53 -233 91
rect -279 19 -273 53
rect -239 19 -233 53
rect -279 -19 -233 19
rect -279 -53 -273 -19
rect -239 -53 -233 -19
rect -279 -91 -233 -53
rect -279 -125 -273 -91
rect -239 -125 -233 -91
rect -279 -163 -233 -125
rect -279 -197 -273 -163
rect -239 -197 -233 -163
rect -279 -235 -233 -197
rect -279 -269 -273 -235
rect -239 -269 -233 -235
rect -279 -307 -233 -269
rect -279 -341 -273 -307
rect -239 -341 -233 -307
rect -279 -386 -233 -341
rect -151 269 -105 314
rect -151 235 -145 269
rect -111 235 -105 269
rect -151 197 -105 235
rect -151 163 -145 197
rect -111 163 -105 197
rect -151 125 -105 163
rect -151 91 -145 125
rect -111 91 -105 125
rect -151 53 -105 91
rect -151 19 -145 53
rect -111 19 -105 53
rect -151 -19 -105 19
rect -151 -53 -145 -19
rect -111 -53 -105 -19
rect -151 -91 -105 -53
rect -151 -125 -145 -91
rect -111 -125 -105 -91
rect -151 -163 -105 -125
rect -151 -197 -145 -163
rect -111 -197 -105 -163
rect -151 -235 -105 -197
rect -151 -269 -145 -235
rect -111 -269 -105 -235
rect -151 -307 -105 -269
rect -151 -341 -145 -307
rect -111 -341 -105 -307
rect -151 -386 -105 -341
rect -23 269 23 314
rect -23 235 -17 269
rect 17 235 23 269
rect -23 197 23 235
rect -23 163 -17 197
rect 17 163 23 197
rect -23 125 23 163
rect -23 91 -17 125
rect 17 91 23 125
rect -23 53 23 91
rect -23 19 -17 53
rect 17 19 23 53
rect -23 -19 23 19
rect -23 -53 -17 -19
rect 17 -53 23 -19
rect -23 -91 23 -53
rect -23 -125 -17 -91
rect 17 -125 23 -91
rect -23 -163 23 -125
rect -23 -197 -17 -163
rect 17 -197 23 -163
rect -23 -235 23 -197
rect -23 -269 -17 -235
rect 17 -269 23 -235
rect -23 -307 23 -269
rect -23 -341 -17 -307
rect 17 -341 23 -307
rect -23 -386 23 -341
rect 105 269 151 314
rect 105 235 111 269
rect 145 235 151 269
rect 105 197 151 235
rect 105 163 111 197
rect 145 163 151 197
rect 105 125 151 163
rect 105 91 111 125
rect 145 91 151 125
rect 105 53 151 91
rect 105 19 111 53
rect 145 19 151 53
rect 105 -19 151 19
rect 105 -53 111 -19
rect 145 -53 151 -19
rect 105 -91 151 -53
rect 105 -125 111 -91
rect 145 -125 151 -91
rect 105 -163 151 -125
rect 105 -197 111 -163
rect 145 -197 151 -163
rect 105 -235 151 -197
rect 105 -269 111 -235
rect 145 -269 151 -235
rect 105 -307 151 -269
rect 105 -341 111 -307
rect 145 -341 151 -307
rect 105 -386 151 -341
rect 233 269 279 314
rect 233 235 239 269
rect 273 235 279 269
rect 233 197 279 235
rect 233 163 239 197
rect 273 163 279 197
rect 233 125 279 163
rect 233 91 239 125
rect 273 91 279 125
rect 233 53 279 91
rect 233 19 239 53
rect 273 19 279 53
rect 233 -19 279 19
rect 233 -53 239 -19
rect 273 -53 279 -19
rect 233 -91 279 -53
rect 233 -125 239 -91
rect 273 -125 279 -91
rect 233 -163 279 -125
rect 233 -197 239 -163
rect 273 -197 279 -163
rect 233 -235 279 -197
rect 233 -269 239 -235
rect 273 -269 279 -235
rect 233 -307 279 -269
rect 233 -341 239 -307
rect 273 -341 279 -307
rect 233 -386 279 -341
rect 361 269 407 314
rect 361 235 367 269
rect 401 235 407 269
rect 361 197 407 235
rect 361 163 367 197
rect 401 163 407 197
rect 361 125 407 163
rect 361 91 367 125
rect 401 91 407 125
rect 361 53 407 91
rect 361 19 367 53
rect 401 19 407 53
rect 361 -19 407 19
rect 361 -53 367 -19
rect 401 -53 407 -19
rect 361 -91 407 -53
rect 361 -125 367 -91
rect 401 -125 407 -91
rect 361 -163 407 -125
rect 361 -197 367 -163
rect 401 -197 407 -163
rect 361 -235 407 -197
rect 361 -269 367 -235
rect 401 -269 407 -235
rect 361 -307 407 -269
rect 361 -341 367 -307
rect 401 -341 407 -307
rect 361 -386 407 -341
rect 489 269 535 314
rect 489 235 495 269
rect 529 235 535 269
rect 489 197 535 235
rect 489 163 495 197
rect 529 163 535 197
rect 489 125 535 163
rect 489 91 495 125
rect 529 91 535 125
rect 489 53 535 91
rect 489 19 495 53
rect 529 19 535 53
rect 489 -19 535 19
rect 489 -53 495 -19
rect 529 -53 535 -19
rect 489 -91 535 -53
rect 489 -125 495 -91
rect 529 -125 535 -91
rect 489 -163 535 -125
rect 489 -197 495 -163
rect 529 -197 535 -163
rect 489 -235 535 -197
rect 489 -269 495 -235
rect 529 -269 535 -235
rect 489 -307 535 -269
rect 489 -341 495 -307
rect 529 -341 535 -307
rect 489 -386 535 -341
rect 617 269 663 314
rect 617 235 623 269
rect 657 235 663 269
rect 617 197 663 235
rect 617 163 623 197
rect 657 163 663 197
rect 617 125 663 163
rect 617 91 623 125
rect 657 91 663 125
rect 617 53 663 91
rect 617 19 623 53
rect 657 19 663 53
rect 617 -19 663 19
rect 617 -53 623 -19
rect 657 -53 663 -19
rect 617 -91 663 -53
rect 617 -125 623 -91
rect 657 -125 663 -91
rect 617 -163 663 -125
rect 617 -197 623 -163
rect 657 -197 663 -163
rect 617 -235 663 -197
rect 617 -269 623 -235
rect 657 -269 663 -235
rect 617 -307 663 -269
rect 617 -341 623 -307
rect 657 -341 663 -307
rect 617 -386 663 -341
rect 745 269 791 314
rect 745 235 751 269
rect 785 235 791 269
rect 745 197 791 235
rect 745 163 751 197
rect 785 163 791 197
rect 745 125 791 163
rect 745 91 751 125
rect 785 91 791 125
rect 745 53 791 91
rect 745 19 751 53
rect 785 19 791 53
rect 745 -19 791 19
rect 745 -53 751 -19
rect 785 -53 791 -19
rect 745 -91 791 -53
rect 745 -125 751 -91
rect 785 -125 791 -91
rect 745 -163 791 -125
rect 745 -197 751 -163
rect 785 -197 791 -163
rect 745 -235 791 -197
rect 745 -269 751 -235
rect 785 -269 791 -235
rect 745 -307 791 -269
rect 745 -341 751 -307
rect 785 -341 791 -307
rect 745 -386 791 -341
rect 873 269 919 314
rect 873 235 879 269
rect 913 235 919 269
rect 873 197 919 235
rect 873 163 879 197
rect 913 163 919 197
rect 873 125 919 163
rect 873 91 879 125
rect 913 91 919 125
rect 873 53 919 91
rect 873 19 879 53
rect 913 19 919 53
rect 873 -19 919 19
rect 873 -53 879 -19
rect 913 -53 919 -19
rect 873 -91 919 -53
rect 873 -125 879 -91
rect 913 -125 919 -91
rect 873 -163 919 -125
rect 873 -197 879 -163
rect 913 -197 919 -163
rect 873 -235 919 -197
rect 873 -269 879 -235
rect 913 -269 919 -235
rect 873 -307 919 -269
rect 873 -341 879 -307
rect 913 -341 919 -307
rect 873 -386 919 -341
rect 1001 269 1047 314
rect 1001 235 1007 269
rect 1041 235 1047 269
rect 1001 197 1047 235
rect 1001 163 1007 197
rect 1041 163 1047 197
rect 1001 125 1047 163
rect 1001 91 1007 125
rect 1041 91 1047 125
rect 1001 53 1047 91
rect 1001 19 1007 53
rect 1041 19 1047 53
rect 1001 -19 1047 19
rect 1001 -53 1007 -19
rect 1041 -53 1047 -19
rect 1001 -91 1047 -53
rect 1001 -125 1007 -91
rect 1041 -125 1047 -91
rect 1001 -163 1047 -125
rect 1001 -197 1007 -163
rect 1041 -197 1047 -163
rect 1001 -235 1047 -197
rect 1001 -269 1007 -235
rect 1041 -269 1047 -235
rect 1001 -307 1047 -269
rect 1001 -341 1007 -307
rect 1041 -341 1047 -307
rect 1001 -386 1047 -341
rect 1129 269 1175 314
rect 1129 235 1135 269
rect 1169 235 1175 269
rect 1129 197 1175 235
rect 1129 163 1135 197
rect 1169 163 1175 197
rect 1129 125 1175 163
rect 1129 91 1135 125
rect 1169 91 1175 125
rect 1129 53 1175 91
rect 1129 19 1135 53
rect 1169 19 1175 53
rect 1129 -19 1175 19
rect 1129 -53 1135 -19
rect 1169 -53 1175 -19
rect 1129 -91 1175 -53
rect 1129 -125 1135 -91
rect 1169 -125 1175 -91
rect 1129 -163 1175 -125
rect 1129 -197 1135 -163
rect 1169 -197 1175 -163
rect 1129 -235 1175 -197
rect 1129 -269 1135 -235
rect 1169 -269 1175 -235
rect 1129 -307 1175 -269
rect 1129 -341 1135 -307
rect 1169 -341 1175 -307
rect 1129 -386 1175 -341
rect 1257 269 1303 314
rect 1257 235 1263 269
rect 1297 235 1303 269
rect 1257 197 1303 235
rect 1257 163 1263 197
rect 1297 163 1303 197
rect 1257 125 1303 163
rect 1257 91 1263 125
rect 1297 91 1303 125
rect 1257 53 1303 91
rect 1257 19 1263 53
rect 1297 19 1303 53
rect 1257 -19 1303 19
rect 1257 -53 1263 -19
rect 1297 -53 1303 -19
rect 1257 -91 1303 -53
rect 1257 -125 1263 -91
rect 1297 -125 1303 -91
rect 1257 -163 1303 -125
rect 1257 -197 1263 -163
rect 1297 -197 1303 -163
rect 1257 -235 1303 -197
rect 1257 -269 1263 -235
rect 1297 -269 1303 -235
rect 1257 -307 1303 -269
rect 1257 -341 1263 -307
rect 1297 -341 1303 -307
rect 1257 -386 1303 -341
rect 1385 269 1431 314
rect 1385 235 1391 269
rect 1425 235 1431 269
rect 1385 197 1431 235
rect 1385 163 1391 197
rect 1425 163 1431 197
rect 1385 125 1431 163
rect 1385 91 1391 125
rect 1425 91 1431 125
rect 1385 53 1431 91
rect 1385 19 1391 53
rect 1425 19 1431 53
rect 1385 -19 1431 19
rect 1385 -53 1391 -19
rect 1425 -53 1431 -19
rect 1385 -91 1431 -53
rect 1385 -125 1391 -91
rect 1425 -125 1431 -91
rect 1385 -163 1431 -125
rect 1385 -197 1391 -163
rect 1425 -197 1431 -163
rect 1385 -235 1431 -197
rect 1385 -269 1391 -235
rect 1425 -269 1431 -235
rect 1385 -307 1431 -269
rect 1385 -341 1391 -307
rect 1425 -341 1431 -307
rect 1385 -386 1431 -341
rect 1513 269 1559 314
rect 1513 235 1519 269
rect 1553 235 1559 269
rect 1513 197 1559 235
rect 1513 163 1519 197
rect 1553 163 1559 197
rect 1513 125 1559 163
rect 1513 91 1519 125
rect 1553 91 1559 125
rect 1513 53 1559 91
rect 1513 19 1519 53
rect 1553 19 1559 53
rect 1513 -19 1559 19
rect 1513 -53 1519 -19
rect 1553 -53 1559 -19
rect 1513 -91 1559 -53
rect 1513 -125 1519 -91
rect 1553 -125 1559 -91
rect 1513 -163 1559 -125
rect 1513 -197 1519 -163
rect 1553 -197 1559 -163
rect 1513 -235 1559 -197
rect 1513 -269 1519 -235
rect 1553 -269 1559 -235
rect 1513 -307 1559 -269
rect 1513 -341 1519 -307
rect 1553 -341 1559 -307
rect 1513 -386 1559 -341
rect 1641 269 1687 314
rect 1641 235 1647 269
rect 1681 235 1687 269
rect 1641 197 1687 235
rect 1641 163 1647 197
rect 1681 163 1687 197
rect 1641 125 1687 163
rect 1641 91 1647 125
rect 1681 91 1687 125
rect 1641 53 1687 91
rect 1641 19 1647 53
rect 1681 19 1687 53
rect 1641 -19 1687 19
rect 1641 -53 1647 -19
rect 1681 -53 1687 -19
rect 1641 -91 1687 -53
rect 1641 -125 1647 -91
rect 1681 -125 1687 -91
rect 1641 -163 1687 -125
rect 1641 -197 1647 -163
rect 1681 -197 1687 -163
rect 1641 -235 1687 -197
rect 1641 -269 1647 -235
rect 1681 -269 1687 -235
rect 1641 -307 1687 -269
rect 1641 -341 1647 -307
rect 1681 -341 1687 -307
rect 1641 -386 1687 -341
rect 1769 269 1815 314
rect 1769 235 1775 269
rect 1809 235 1815 269
rect 1769 197 1815 235
rect 1769 163 1775 197
rect 1809 163 1815 197
rect 1769 125 1815 163
rect 1769 91 1775 125
rect 1809 91 1815 125
rect 1769 53 1815 91
rect 1769 19 1775 53
rect 1809 19 1815 53
rect 1769 -19 1815 19
rect 1769 -53 1775 -19
rect 1809 -53 1815 -19
rect 1769 -91 1815 -53
rect 1769 -125 1775 -91
rect 1809 -125 1815 -91
rect 1769 -163 1815 -125
rect 1769 -197 1775 -163
rect 1809 -197 1815 -163
rect 1769 -235 1815 -197
rect 1769 -269 1775 -235
rect 1809 -269 1815 -235
rect 1769 -307 1815 -269
rect 1769 -341 1775 -307
rect 1809 -341 1815 -307
rect 1769 -386 1815 -341
rect 1897 269 1943 314
rect 1897 235 1903 269
rect 1937 235 1943 269
rect 1897 197 1943 235
rect 1897 163 1903 197
rect 1937 163 1943 197
rect 1897 125 1943 163
rect 1897 91 1903 125
rect 1937 91 1943 125
rect 1897 53 1943 91
rect 1897 19 1903 53
rect 1937 19 1943 53
rect 1897 -19 1943 19
rect 1897 -53 1903 -19
rect 1937 -53 1943 -19
rect 1897 -91 1943 -53
rect 1897 -125 1903 -91
rect 1937 -125 1943 -91
rect 1897 -163 1943 -125
rect 1897 -197 1903 -163
rect 1937 -197 1943 -163
rect 1897 -235 1943 -197
rect 1897 -269 1903 -235
rect 1937 -269 1943 -235
rect 1897 -307 1943 -269
rect 1897 -341 1903 -307
rect 1937 -341 1943 -307
rect 1897 -386 1943 -341
rect 2025 269 2071 314
rect 2025 235 2031 269
rect 2065 235 2071 269
rect 2025 197 2071 235
rect 2025 163 2031 197
rect 2065 163 2071 197
rect 2025 125 2071 163
rect 2025 91 2031 125
rect 2065 91 2071 125
rect 2025 53 2071 91
rect 2025 19 2031 53
rect 2065 19 2071 53
rect 2025 -19 2071 19
rect 2025 -53 2031 -19
rect 2065 -53 2071 -19
rect 2025 -91 2071 -53
rect 2025 -125 2031 -91
rect 2065 -125 2071 -91
rect 2025 -163 2071 -125
rect 2025 -197 2031 -163
rect 2065 -197 2071 -163
rect 2025 -235 2071 -197
rect 2025 -269 2031 -235
rect 2065 -269 2071 -235
rect 2025 -307 2071 -269
rect 2025 -341 2031 -307
rect 2065 -341 2071 -307
rect 2025 -386 2071 -341
rect 2153 269 2199 314
rect 2153 235 2159 269
rect 2193 235 2199 269
rect 2153 197 2199 235
rect 2153 163 2159 197
rect 2193 163 2199 197
rect 2153 125 2199 163
rect 2153 91 2159 125
rect 2193 91 2199 125
rect 2153 53 2199 91
rect 2153 19 2159 53
rect 2193 19 2199 53
rect 2153 -19 2199 19
rect 2153 -53 2159 -19
rect 2193 -53 2199 -19
rect 2153 -91 2199 -53
rect 2153 -125 2159 -91
rect 2193 -125 2199 -91
rect 2153 -163 2199 -125
rect 2153 -197 2159 -163
rect 2193 -197 2199 -163
rect 2153 -235 2199 -197
rect 2153 -269 2159 -235
rect 2193 -269 2199 -235
rect 2153 -307 2199 -269
rect 2153 -341 2159 -307
rect 2193 -341 2199 -307
rect 2153 -386 2199 -341
rect 2281 269 2327 314
rect 2281 235 2287 269
rect 2321 235 2327 269
rect 2281 197 2327 235
rect 2281 163 2287 197
rect 2321 163 2327 197
rect 2281 125 2327 163
rect 2281 91 2287 125
rect 2321 91 2327 125
rect 2281 53 2327 91
rect 2281 19 2287 53
rect 2321 19 2327 53
rect 2281 -19 2327 19
rect 2281 -53 2287 -19
rect 2321 -53 2327 -19
rect 2281 -91 2327 -53
rect 2281 -125 2287 -91
rect 2321 -125 2327 -91
rect 2281 -163 2327 -125
rect 2281 -197 2287 -163
rect 2321 -197 2327 -163
rect 2281 -235 2327 -197
rect 2281 -269 2287 -235
rect 2321 -269 2327 -235
rect 2281 -307 2327 -269
rect 2281 -341 2287 -307
rect 2321 -341 2327 -307
rect 2281 -386 2327 -341
rect 2409 269 2455 314
rect 2409 235 2415 269
rect 2449 235 2455 269
rect 2409 197 2455 235
rect 2409 163 2415 197
rect 2449 163 2455 197
rect 2409 125 2455 163
rect 2409 91 2415 125
rect 2449 91 2455 125
rect 2409 53 2455 91
rect 2409 19 2415 53
rect 2449 19 2455 53
rect 2409 -19 2455 19
rect 2409 -53 2415 -19
rect 2449 -53 2455 -19
rect 2409 -91 2455 -53
rect 2409 -125 2415 -91
rect 2449 -125 2455 -91
rect 2409 -163 2455 -125
rect 2409 -197 2415 -163
rect 2449 -197 2455 -163
rect 2409 -235 2455 -197
rect 2409 -269 2415 -235
rect 2449 -269 2455 -235
rect 2409 -307 2455 -269
rect 2409 -341 2415 -307
rect 2449 -341 2455 -307
rect 2409 -386 2455 -341
rect 2537 269 2583 314
rect 2537 235 2543 269
rect 2577 235 2583 269
rect 2537 197 2583 235
rect 2537 163 2543 197
rect 2577 163 2583 197
rect 2537 125 2583 163
rect 2537 91 2543 125
rect 2577 91 2583 125
rect 2537 53 2583 91
rect 2537 19 2543 53
rect 2577 19 2583 53
rect 2537 -19 2583 19
rect 2537 -53 2543 -19
rect 2577 -53 2583 -19
rect 2537 -91 2583 -53
rect 2537 -125 2543 -91
rect 2577 -125 2583 -91
rect 2537 -163 2583 -125
rect 2537 -197 2543 -163
rect 2577 -197 2583 -163
rect 2537 -235 2583 -197
rect 2537 -269 2543 -235
rect 2577 -269 2583 -235
rect 2537 -307 2583 -269
rect 2537 -341 2543 -307
rect 2577 -341 2583 -307
rect 2537 -386 2583 -341
<< labels >>
flabel metal1 s -2496 378 -2496 378 0 FreeSans 300 0 0 0 G
port 1 nsew
flabel metal1 s -2368 378 -2368 378 0 FreeSans 300 0 0 0 G
port 1 nsew
flabel metal1 s -2240 378 -2240 378 0 FreeSans 300 0 0 0 G
port 1 nsew
flabel metal1 s -2112 378 -2112 378 0 FreeSans 300 0 0 0 G
port 1 nsew
flabel metal1 s -1984 378 -1984 378 0 FreeSans 300 0 0 0 G
port 1 nsew
flabel metal1 s -1855 378 -1855 378 0 FreeSans 300 0 0 0 G
port 1 nsew
flabel metal1 s -1728 378 -1728 378 0 FreeSans 300 0 0 0 G
port 1 nsew
flabel metal1 s -1600 378 -1600 378 0 FreeSans 300 0 0 0 G
port 1 nsew
flabel metal1 s -1472 378 -1472 378 0 FreeSans 300 0 0 0 G
port 1 nsew
flabel metal1 s -1344 378 -1344 378 0 FreeSans 300 0 0 0 G
port 1 nsew
flabel metal1 s -1216 378 -1216 378 0 FreeSans 300 0 0 0 G
port 1 nsew
flabel metal1 s -1088 378 -1088 378 0 FreeSans 300 0 0 0 G
port 1 nsew
flabel metal1 s -960 378 -960 378 0 FreeSans 300 0 0 0 G
port 1 nsew
flabel metal1 s -832 378 -832 378 0 FreeSans 300 0 0 0 G
port 1 nsew
flabel metal1 s -704 378 -704 378 0 FreeSans 300 0 0 0 G
port 1 nsew
flabel metal1 s -576 378 -576 378 0 FreeSans 300 0 0 0 G
port 1 nsew
flabel metal1 s -448 378 -448 378 0 FreeSans 300 0 0 0 G
port 1 nsew
flabel metal1 s -320 378 -320 378 0 FreeSans 300 0 0 0 G
port 1 nsew
flabel metal1 s -192 378 -192 378 0 FreeSans 300 0 0 0 G
port 1 nsew
flabel metal1 s -64 378 -64 378 0 FreeSans 300 0 0 0 G
port 1 nsew
flabel metal1 s 64 378 64 378 0 FreeSans 300 0 0 0 G
port 1 nsew
flabel metal1 s 192 378 192 378 0 FreeSans 300 0 0 0 G
port 1 nsew
flabel metal1 s 320 378 320 378 0 FreeSans 300 0 0 0 G
port 1 nsew
flabel metal1 s 448 378 448 378 0 FreeSans 300 0 0 0 G
port 1 nsew
flabel metal1 s 576 378 576 378 0 FreeSans 300 0 0 0 G
port 1 nsew
flabel metal1 s 704 378 704 378 0 FreeSans 300 0 0 0 G
port 1 nsew
flabel metal1 s 832 378 832 378 0 FreeSans 300 0 0 0 G
port 1 nsew
flabel metal1 s 960 378 960 378 0 FreeSans 300 0 0 0 G
port 1 nsew
flabel metal1 s 1088 378 1088 378 0 FreeSans 300 0 0 0 G
port 1 nsew
flabel metal1 s 1216 378 1216 378 0 FreeSans 300 0 0 0 G
port 1 nsew
flabel metal1 s 1344 378 1344 378 0 FreeSans 300 0 0 0 G
port 1 nsew
flabel metal1 s 1472 378 1472 378 0 FreeSans 300 0 0 0 G
port 1 nsew
flabel metal1 s 1600 378 1600 378 0 FreeSans 300 0 0 0 G
port 1 nsew
flabel metal1 s 1728 378 1728 378 0 FreeSans 300 0 0 0 G
port 1 nsew
flabel metal1 s 1855 378 1855 378 0 FreeSans 300 0 0 0 G
port 1 nsew
flabel metal1 s 1984 378 1984 378 0 FreeSans 300 0 0 0 G
port 1 nsew
flabel metal1 s 2112 378 2112 378 0 FreeSans 300 0 0 0 G
port 1 nsew
flabel metal1 s 2240 378 2240 378 0 FreeSans 300 0 0 0 G
port 1 nsew
flabel metal1 s 2368 378 2368 378 0 FreeSans 300 0 0 0 G
port 1 nsew
flabel metal1 s 2496 378 2496 378 0 FreeSans 300 0 0 0 G
port 1 nsew
flabel metal1 s -2560 -36 -2560 -36 0 FreeSans 300 0 0 0 D
port 2 nsew
flabel metal1 s -2432 -36 -2432 -36 0 FreeSans 300 0 0 0 S
port 3 nsew
flabel metal1 s -2304 -36 -2304 -36 0 FreeSans 300 0 0 0 D
port 2 nsew
flabel metal1 s -2176 -36 -2176 -36 0 FreeSans 300 0 0 0 S
port 3 nsew
flabel metal1 s -2048 -36 -2048 -36 0 FreeSans 300 0 0 0 D
port 2 nsew
flabel metal1 s -1920 -36 -1920 -36 0 FreeSans 300 0 0 0 S
port 3 nsew
flabel metal1 s -1792 -36 -1792 -36 0 FreeSans 300 0 0 0 D
port 2 nsew
flabel metal1 s -1664 -36 -1664 -36 0 FreeSans 300 0 0 0 S
port 3 nsew
flabel metal1 s -1536 -36 -1536 -36 0 FreeSans 300 0 0 0 D
port 2 nsew
flabel metal1 s -1408 -36 -1408 -36 0 FreeSans 300 0 0 0 S
port 3 nsew
flabel metal1 s -1280 -36 -1280 -36 0 FreeSans 300 0 0 0 D
port 2 nsew
flabel metal1 s -1152 -36 -1152 -36 0 FreeSans 300 0 0 0 S
port 3 nsew
flabel metal1 s -1024 -36 -1024 -36 0 FreeSans 300 0 0 0 D
port 2 nsew
flabel metal1 s -896 -36 -896 -36 0 FreeSans 300 0 0 0 S
port 3 nsew
flabel metal1 s -768 -36 -768 -36 0 FreeSans 300 0 0 0 D
port 2 nsew
flabel metal1 s -640 -36 -640 -36 0 FreeSans 300 0 0 0 S
port 3 nsew
flabel metal1 s -512 -36 -512 -36 0 FreeSans 300 0 0 0 D
port 2 nsew
flabel metal1 s -384 -36 -384 -36 0 FreeSans 300 0 0 0 S
port 3 nsew
flabel metal1 s -256 -36 -256 -36 0 FreeSans 300 0 0 0 D
port 2 nsew
flabel metal1 s -128 -36 -128 -36 0 FreeSans 300 0 0 0 S
port 3 nsew
flabel metal1 s 0 -36 0 -36 0 FreeSans 300 0 0 0 D
port 2 nsew
flabel metal1 s 128 -36 128 -36 0 FreeSans 300 0 0 0 S
port 3 nsew
flabel metal1 s 256 -36 256 -36 0 FreeSans 300 0 0 0 D
port 2 nsew
flabel metal1 s 384 -36 384 -36 0 FreeSans 300 0 0 0 S
port 3 nsew
flabel metal1 s 512 -36 512 -36 0 FreeSans 300 0 0 0 D
port 2 nsew
flabel metal1 s 640 -36 640 -36 0 FreeSans 300 0 0 0 S
port 3 nsew
flabel metal1 s 768 -36 768 -36 0 FreeSans 300 0 0 0 D
port 2 nsew
flabel metal1 s 896 -36 896 -36 0 FreeSans 300 0 0 0 S
port 3 nsew
flabel metal1 s 1024 -36 1024 -36 0 FreeSans 300 0 0 0 D
port 2 nsew
flabel metal1 s 1152 -36 1152 -36 0 FreeSans 300 0 0 0 S
port 3 nsew
flabel metal1 s 1280 -36 1280 -36 0 FreeSans 300 0 0 0 D
port 2 nsew
flabel metal1 s 1408 -36 1408 -36 0 FreeSans 300 0 0 0 S
port 3 nsew
flabel metal1 s 1536 -36 1536 -36 0 FreeSans 300 0 0 0 D
port 2 nsew
flabel metal1 s 1664 -36 1664 -36 0 FreeSans 300 0 0 0 S
port 3 nsew
flabel metal1 s 1792 -36 1792 -36 0 FreeSans 300 0 0 0 D
port 2 nsew
flabel metal1 s 1920 -36 1920 -36 0 FreeSans 300 0 0 0 S
port 3 nsew
flabel metal1 s 2048 -36 2048 -36 0 FreeSans 300 0 0 0 D
port 2 nsew
flabel metal1 s 2176 -36 2176 -36 0 FreeSans 300 0 0 0 S
port 3 nsew
flabel metal1 s 2304 -36 2304 -36 0 FreeSans 300 0 0 0 D
port 2 nsew
flabel metal1 s 2432 -36 2432 -36 0 FreeSans 300 0 0 0 S
port 3 nsew
flabel metal1 s 2560 -36 2560 -36 0 FreeSans 300 0 0 0 D
port 2 nsew
<< properties >>
string FIXED_BBOX -2674 -481 2674 481
<< end >>
