magic
tech sky130A
magscale 1 2
timestamp 1679988683
<< checkpaint >>
rect -1518 -2321 1518 2321
<< pwell >>
rect -258 -1061 258 1061
<< ndiff >>
rect -100 891 100 903
rect -100 857 -88 891
rect 88 857 100 891
rect -100 800 100 857
rect -100 -857 100 -800
rect -100 -891 -88 -857
rect 88 -891 100 -857
rect -100 -903 100 -891
<< ndiffc >>
rect -88 857 88 891
rect -88 -891 88 -857
<< psubdiff >>
rect -222 991 -126 1025
rect 126 991 222 1025
rect -222 929 -188 991
rect 188 929 222 991
rect -222 -991 -188 -929
rect 188 -991 222 -929
rect -222 -1025 -126 -991
rect 126 -1025 222 -991
<< psubdiffcont >>
rect -126 991 126 1025
rect -222 -929 -188 929
rect 188 -929 222 929
rect -126 -1025 126 -991
<< ndiffres >>
rect -100 -800 100 800
<< locali >>
rect -222 991 -126 1025
rect 126 991 222 1025
rect -222 929 -188 991
rect 188 929 222 991
rect -104 857 -88 891
rect 88 857 104 891
rect -104 -891 -88 -857
rect 88 -891 104 -857
rect -222 -991 -188 -929
rect 188 -991 222 -929
rect -222 -1025 -126 -991
rect 126 -1025 222 -991
<< viali >>
rect -88 857 88 891
rect -88 817 88 857
rect -88 -857 88 -817
rect -88 -891 88 -857
<< metal1 >>
rect -100 891 100 897
rect -100 817 -88 891
rect 88 817 100 891
rect -100 811 100 817
rect -100 -817 100 -811
rect -100 -891 -88 -817
rect 88 -891 100 -817
rect -100 -897 100 -891
<< labels >>
flabel metal1 0 853 0 853 0 FreeSans 240 0 0 0 1
flabel metal1 0 -853 0 -853 0 FreeSans 240 0 0 0 2
<< properties >>
string FIXED_BBOX -205 -1008 205 1008
<< end >>

