magic
tech sky130A
magscale 1 2
timestamp 1680002671
<< error_p >>
rect -2015 391 -1953 397
rect -1887 391 -1825 397
rect -1759 391 -1697 397
rect -1631 391 -1569 397
rect -1503 391 -1441 397
rect -1375 391 -1313 397
rect -1247 391 -1185 397
rect -1119 391 -1057 397
rect -991 391 -929 397
rect -863 391 -801 397
rect -735 391 -673 397
rect -607 391 -545 397
rect -479 391 -417 397
rect -351 391 -289 397
rect -223 391 -161 397
rect -95 391 -33 397
rect 33 391 95 397
rect 161 391 223 397
rect 289 391 351 397
rect 417 391 479 397
rect 545 391 607 397
rect 673 391 735 397
rect 801 391 863 397
rect 929 391 991 397
rect 1057 391 1119 397
rect 1185 391 1247 397
rect 1313 391 1375 397
rect 1441 391 1503 397
rect 1569 391 1631 397
rect 1697 391 1759 397
rect 1825 391 1887 397
rect 1953 391 2015 397
rect -2015 357 -2001 391
rect -1887 357 -1873 391
rect -1759 357 -1745 391
rect -1631 357 -1617 391
rect -1503 357 -1489 391
rect -1375 357 -1361 391
rect -1247 357 -1233 391
rect -1119 357 -1105 391
rect -991 357 -977 391
rect -863 357 -849 391
rect -735 357 -721 391
rect -607 357 -593 391
rect -479 357 -465 391
rect -351 357 -337 391
rect -223 357 -209 391
rect -95 357 -81 391
rect 33 357 47 391
rect 161 357 175 391
rect 289 357 303 391
rect 417 357 431 391
rect 545 357 559 391
rect 673 357 687 391
rect 801 357 815 391
rect 929 357 943 391
rect 1057 357 1071 391
rect 1185 357 1199 391
rect 1313 357 1327 391
rect 1441 357 1455 391
rect 1569 357 1583 391
rect 1697 357 1711 391
rect 1825 357 1839 391
rect 1953 357 1967 391
rect -2015 351 -1953 357
rect -1887 351 -1825 357
rect -1759 351 -1697 357
rect -1631 351 -1569 357
rect -1503 351 -1441 357
rect -1375 351 -1313 357
rect -1247 351 -1185 357
rect -1119 351 -1057 357
rect -991 351 -929 357
rect -863 351 -801 357
rect -735 351 -673 357
rect -607 351 -545 357
rect -479 351 -417 357
rect -351 351 -289 357
rect -223 351 -161 357
rect -95 351 -33 357
rect 33 351 95 357
rect 161 351 223 357
rect 289 351 351 357
rect 417 351 479 357
rect 545 351 607 357
rect 673 351 735 357
rect 801 351 863 357
rect 929 351 991 357
rect 1057 351 1119 357
rect 1185 351 1247 357
rect 1313 351 1375 357
rect 1441 351 1503 357
rect 1569 351 1631 357
rect 1697 351 1759 357
rect 1825 351 1887 357
rect 1953 351 2015 357
<< pwell >>
rect -2205 -519 2205 519
<< nmoslvt >>
rect -2019 -381 -1949 319
rect -1891 -381 -1821 319
rect -1763 -381 -1693 319
rect -1635 -381 -1565 319
rect -1507 -381 -1437 319
rect -1379 -381 -1309 319
rect -1251 -381 -1181 319
rect -1123 -381 -1053 319
rect -995 -381 -925 319
rect -867 -381 -797 319
rect -739 -381 -669 319
rect -611 -381 -541 319
rect -483 -381 -413 319
rect -355 -381 -285 319
rect -227 -381 -157 319
rect -99 -381 -29 319
rect 29 -381 99 319
rect 157 -381 227 319
rect 285 -381 355 319
rect 413 -381 483 319
rect 541 -381 611 319
rect 669 -381 739 319
rect 797 -381 867 319
rect 925 -381 995 319
rect 1053 -381 1123 319
rect 1181 -381 1251 319
rect 1309 -381 1379 319
rect 1437 -381 1507 319
rect 1565 -381 1635 319
rect 1693 -381 1763 319
rect 1821 -381 1891 319
rect 1949 -381 2019 319
<< ndiff >>
rect -2077 292 -2019 319
rect -2077 258 -2065 292
rect -2031 258 -2019 292
rect -2077 224 -2019 258
rect -2077 190 -2065 224
rect -2031 190 -2019 224
rect -2077 156 -2019 190
rect -2077 122 -2065 156
rect -2031 122 -2019 156
rect -2077 88 -2019 122
rect -2077 54 -2065 88
rect -2031 54 -2019 88
rect -2077 20 -2019 54
rect -2077 -14 -2065 20
rect -2031 -14 -2019 20
rect -2077 -48 -2019 -14
rect -2077 -82 -2065 -48
rect -2031 -82 -2019 -48
rect -2077 -116 -2019 -82
rect -2077 -150 -2065 -116
rect -2031 -150 -2019 -116
rect -2077 -184 -2019 -150
rect -2077 -218 -2065 -184
rect -2031 -218 -2019 -184
rect -2077 -252 -2019 -218
rect -2077 -286 -2065 -252
rect -2031 -286 -2019 -252
rect -2077 -320 -2019 -286
rect -2077 -354 -2065 -320
rect -2031 -354 -2019 -320
rect -2077 -381 -2019 -354
rect -1949 292 -1891 319
rect -1949 258 -1937 292
rect -1903 258 -1891 292
rect -1949 224 -1891 258
rect -1949 190 -1937 224
rect -1903 190 -1891 224
rect -1949 156 -1891 190
rect -1949 122 -1937 156
rect -1903 122 -1891 156
rect -1949 88 -1891 122
rect -1949 54 -1937 88
rect -1903 54 -1891 88
rect -1949 20 -1891 54
rect -1949 -14 -1937 20
rect -1903 -14 -1891 20
rect -1949 -48 -1891 -14
rect -1949 -82 -1937 -48
rect -1903 -82 -1891 -48
rect -1949 -116 -1891 -82
rect -1949 -150 -1937 -116
rect -1903 -150 -1891 -116
rect -1949 -184 -1891 -150
rect -1949 -218 -1937 -184
rect -1903 -218 -1891 -184
rect -1949 -252 -1891 -218
rect -1949 -286 -1937 -252
rect -1903 -286 -1891 -252
rect -1949 -320 -1891 -286
rect -1949 -354 -1937 -320
rect -1903 -354 -1891 -320
rect -1949 -381 -1891 -354
rect -1821 292 -1763 319
rect -1821 258 -1809 292
rect -1775 258 -1763 292
rect -1821 224 -1763 258
rect -1821 190 -1809 224
rect -1775 190 -1763 224
rect -1821 156 -1763 190
rect -1821 122 -1809 156
rect -1775 122 -1763 156
rect -1821 88 -1763 122
rect -1821 54 -1809 88
rect -1775 54 -1763 88
rect -1821 20 -1763 54
rect -1821 -14 -1809 20
rect -1775 -14 -1763 20
rect -1821 -48 -1763 -14
rect -1821 -82 -1809 -48
rect -1775 -82 -1763 -48
rect -1821 -116 -1763 -82
rect -1821 -150 -1809 -116
rect -1775 -150 -1763 -116
rect -1821 -184 -1763 -150
rect -1821 -218 -1809 -184
rect -1775 -218 -1763 -184
rect -1821 -252 -1763 -218
rect -1821 -286 -1809 -252
rect -1775 -286 -1763 -252
rect -1821 -320 -1763 -286
rect -1821 -354 -1809 -320
rect -1775 -354 -1763 -320
rect -1821 -381 -1763 -354
rect -1693 292 -1635 319
rect -1693 258 -1681 292
rect -1647 258 -1635 292
rect -1693 224 -1635 258
rect -1693 190 -1681 224
rect -1647 190 -1635 224
rect -1693 156 -1635 190
rect -1693 122 -1681 156
rect -1647 122 -1635 156
rect -1693 88 -1635 122
rect -1693 54 -1681 88
rect -1647 54 -1635 88
rect -1693 20 -1635 54
rect -1693 -14 -1681 20
rect -1647 -14 -1635 20
rect -1693 -48 -1635 -14
rect -1693 -82 -1681 -48
rect -1647 -82 -1635 -48
rect -1693 -116 -1635 -82
rect -1693 -150 -1681 -116
rect -1647 -150 -1635 -116
rect -1693 -184 -1635 -150
rect -1693 -218 -1681 -184
rect -1647 -218 -1635 -184
rect -1693 -252 -1635 -218
rect -1693 -286 -1681 -252
rect -1647 -286 -1635 -252
rect -1693 -320 -1635 -286
rect -1693 -354 -1681 -320
rect -1647 -354 -1635 -320
rect -1693 -381 -1635 -354
rect -1565 292 -1507 319
rect -1565 258 -1553 292
rect -1519 258 -1507 292
rect -1565 224 -1507 258
rect -1565 190 -1553 224
rect -1519 190 -1507 224
rect -1565 156 -1507 190
rect -1565 122 -1553 156
rect -1519 122 -1507 156
rect -1565 88 -1507 122
rect -1565 54 -1553 88
rect -1519 54 -1507 88
rect -1565 20 -1507 54
rect -1565 -14 -1553 20
rect -1519 -14 -1507 20
rect -1565 -48 -1507 -14
rect -1565 -82 -1553 -48
rect -1519 -82 -1507 -48
rect -1565 -116 -1507 -82
rect -1565 -150 -1553 -116
rect -1519 -150 -1507 -116
rect -1565 -184 -1507 -150
rect -1565 -218 -1553 -184
rect -1519 -218 -1507 -184
rect -1565 -252 -1507 -218
rect -1565 -286 -1553 -252
rect -1519 -286 -1507 -252
rect -1565 -320 -1507 -286
rect -1565 -354 -1553 -320
rect -1519 -354 -1507 -320
rect -1565 -381 -1507 -354
rect -1437 292 -1379 319
rect -1437 258 -1425 292
rect -1391 258 -1379 292
rect -1437 224 -1379 258
rect -1437 190 -1425 224
rect -1391 190 -1379 224
rect -1437 156 -1379 190
rect -1437 122 -1425 156
rect -1391 122 -1379 156
rect -1437 88 -1379 122
rect -1437 54 -1425 88
rect -1391 54 -1379 88
rect -1437 20 -1379 54
rect -1437 -14 -1425 20
rect -1391 -14 -1379 20
rect -1437 -48 -1379 -14
rect -1437 -82 -1425 -48
rect -1391 -82 -1379 -48
rect -1437 -116 -1379 -82
rect -1437 -150 -1425 -116
rect -1391 -150 -1379 -116
rect -1437 -184 -1379 -150
rect -1437 -218 -1425 -184
rect -1391 -218 -1379 -184
rect -1437 -252 -1379 -218
rect -1437 -286 -1425 -252
rect -1391 -286 -1379 -252
rect -1437 -320 -1379 -286
rect -1437 -354 -1425 -320
rect -1391 -354 -1379 -320
rect -1437 -381 -1379 -354
rect -1309 292 -1251 319
rect -1309 258 -1297 292
rect -1263 258 -1251 292
rect -1309 224 -1251 258
rect -1309 190 -1297 224
rect -1263 190 -1251 224
rect -1309 156 -1251 190
rect -1309 122 -1297 156
rect -1263 122 -1251 156
rect -1309 88 -1251 122
rect -1309 54 -1297 88
rect -1263 54 -1251 88
rect -1309 20 -1251 54
rect -1309 -14 -1297 20
rect -1263 -14 -1251 20
rect -1309 -48 -1251 -14
rect -1309 -82 -1297 -48
rect -1263 -82 -1251 -48
rect -1309 -116 -1251 -82
rect -1309 -150 -1297 -116
rect -1263 -150 -1251 -116
rect -1309 -184 -1251 -150
rect -1309 -218 -1297 -184
rect -1263 -218 -1251 -184
rect -1309 -252 -1251 -218
rect -1309 -286 -1297 -252
rect -1263 -286 -1251 -252
rect -1309 -320 -1251 -286
rect -1309 -354 -1297 -320
rect -1263 -354 -1251 -320
rect -1309 -381 -1251 -354
rect -1181 292 -1123 319
rect -1181 258 -1169 292
rect -1135 258 -1123 292
rect -1181 224 -1123 258
rect -1181 190 -1169 224
rect -1135 190 -1123 224
rect -1181 156 -1123 190
rect -1181 122 -1169 156
rect -1135 122 -1123 156
rect -1181 88 -1123 122
rect -1181 54 -1169 88
rect -1135 54 -1123 88
rect -1181 20 -1123 54
rect -1181 -14 -1169 20
rect -1135 -14 -1123 20
rect -1181 -48 -1123 -14
rect -1181 -82 -1169 -48
rect -1135 -82 -1123 -48
rect -1181 -116 -1123 -82
rect -1181 -150 -1169 -116
rect -1135 -150 -1123 -116
rect -1181 -184 -1123 -150
rect -1181 -218 -1169 -184
rect -1135 -218 -1123 -184
rect -1181 -252 -1123 -218
rect -1181 -286 -1169 -252
rect -1135 -286 -1123 -252
rect -1181 -320 -1123 -286
rect -1181 -354 -1169 -320
rect -1135 -354 -1123 -320
rect -1181 -381 -1123 -354
rect -1053 292 -995 319
rect -1053 258 -1041 292
rect -1007 258 -995 292
rect -1053 224 -995 258
rect -1053 190 -1041 224
rect -1007 190 -995 224
rect -1053 156 -995 190
rect -1053 122 -1041 156
rect -1007 122 -995 156
rect -1053 88 -995 122
rect -1053 54 -1041 88
rect -1007 54 -995 88
rect -1053 20 -995 54
rect -1053 -14 -1041 20
rect -1007 -14 -995 20
rect -1053 -48 -995 -14
rect -1053 -82 -1041 -48
rect -1007 -82 -995 -48
rect -1053 -116 -995 -82
rect -1053 -150 -1041 -116
rect -1007 -150 -995 -116
rect -1053 -184 -995 -150
rect -1053 -218 -1041 -184
rect -1007 -218 -995 -184
rect -1053 -252 -995 -218
rect -1053 -286 -1041 -252
rect -1007 -286 -995 -252
rect -1053 -320 -995 -286
rect -1053 -354 -1041 -320
rect -1007 -354 -995 -320
rect -1053 -381 -995 -354
rect -925 292 -867 319
rect -925 258 -913 292
rect -879 258 -867 292
rect -925 224 -867 258
rect -925 190 -913 224
rect -879 190 -867 224
rect -925 156 -867 190
rect -925 122 -913 156
rect -879 122 -867 156
rect -925 88 -867 122
rect -925 54 -913 88
rect -879 54 -867 88
rect -925 20 -867 54
rect -925 -14 -913 20
rect -879 -14 -867 20
rect -925 -48 -867 -14
rect -925 -82 -913 -48
rect -879 -82 -867 -48
rect -925 -116 -867 -82
rect -925 -150 -913 -116
rect -879 -150 -867 -116
rect -925 -184 -867 -150
rect -925 -218 -913 -184
rect -879 -218 -867 -184
rect -925 -252 -867 -218
rect -925 -286 -913 -252
rect -879 -286 -867 -252
rect -925 -320 -867 -286
rect -925 -354 -913 -320
rect -879 -354 -867 -320
rect -925 -381 -867 -354
rect -797 292 -739 319
rect -797 258 -785 292
rect -751 258 -739 292
rect -797 224 -739 258
rect -797 190 -785 224
rect -751 190 -739 224
rect -797 156 -739 190
rect -797 122 -785 156
rect -751 122 -739 156
rect -797 88 -739 122
rect -797 54 -785 88
rect -751 54 -739 88
rect -797 20 -739 54
rect -797 -14 -785 20
rect -751 -14 -739 20
rect -797 -48 -739 -14
rect -797 -82 -785 -48
rect -751 -82 -739 -48
rect -797 -116 -739 -82
rect -797 -150 -785 -116
rect -751 -150 -739 -116
rect -797 -184 -739 -150
rect -797 -218 -785 -184
rect -751 -218 -739 -184
rect -797 -252 -739 -218
rect -797 -286 -785 -252
rect -751 -286 -739 -252
rect -797 -320 -739 -286
rect -797 -354 -785 -320
rect -751 -354 -739 -320
rect -797 -381 -739 -354
rect -669 292 -611 319
rect -669 258 -657 292
rect -623 258 -611 292
rect -669 224 -611 258
rect -669 190 -657 224
rect -623 190 -611 224
rect -669 156 -611 190
rect -669 122 -657 156
rect -623 122 -611 156
rect -669 88 -611 122
rect -669 54 -657 88
rect -623 54 -611 88
rect -669 20 -611 54
rect -669 -14 -657 20
rect -623 -14 -611 20
rect -669 -48 -611 -14
rect -669 -82 -657 -48
rect -623 -82 -611 -48
rect -669 -116 -611 -82
rect -669 -150 -657 -116
rect -623 -150 -611 -116
rect -669 -184 -611 -150
rect -669 -218 -657 -184
rect -623 -218 -611 -184
rect -669 -252 -611 -218
rect -669 -286 -657 -252
rect -623 -286 -611 -252
rect -669 -320 -611 -286
rect -669 -354 -657 -320
rect -623 -354 -611 -320
rect -669 -381 -611 -354
rect -541 292 -483 319
rect -541 258 -529 292
rect -495 258 -483 292
rect -541 224 -483 258
rect -541 190 -529 224
rect -495 190 -483 224
rect -541 156 -483 190
rect -541 122 -529 156
rect -495 122 -483 156
rect -541 88 -483 122
rect -541 54 -529 88
rect -495 54 -483 88
rect -541 20 -483 54
rect -541 -14 -529 20
rect -495 -14 -483 20
rect -541 -48 -483 -14
rect -541 -82 -529 -48
rect -495 -82 -483 -48
rect -541 -116 -483 -82
rect -541 -150 -529 -116
rect -495 -150 -483 -116
rect -541 -184 -483 -150
rect -541 -218 -529 -184
rect -495 -218 -483 -184
rect -541 -252 -483 -218
rect -541 -286 -529 -252
rect -495 -286 -483 -252
rect -541 -320 -483 -286
rect -541 -354 -529 -320
rect -495 -354 -483 -320
rect -541 -381 -483 -354
rect -413 292 -355 319
rect -413 258 -401 292
rect -367 258 -355 292
rect -413 224 -355 258
rect -413 190 -401 224
rect -367 190 -355 224
rect -413 156 -355 190
rect -413 122 -401 156
rect -367 122 -355 156
rect -413 88 -355 122
rect -413 54 -401 88
rect -367 54 -355 88
rect -413 20 -355 54
rect -413 -14 -401 20
rect -367 -14 -355 20
rect -413 -48 -355 -14
rect -413 -82 -401 -48
rect -367 -82 -355 -48
rect -413 -116 -355 -82
rect -413 -150 -401 -116
rect -367 -150 -355 -116
rect -413 -184 -355 -150
rect -413 -218 -401 -184
rect -367 -218 -355 -184
rect -413 -252 -355 -218
rect -413 -286 -401 -252
rect -367 -286 -355 -252
rect -413 -320 -355 -286
rect -413 -354 -401 -320
rect -367 -354 -355 -320
rect -413 -381 -355 -354
rect -285 292 -227 319
rect -285 258 -273 292
rect -239 258 -227 292
rect -285 224 -227 258
rect -285 190 -273 224
rect -239 190 -227 224
rect -285 156 -227 190
rect -285 122 -273 156
rect -239 122 -227 156
rect -285 88 -227 122
rect -285 54 -273 88
rect -239 54 -227 88
rect -285 20 -227 54
rect -285 -14 -273 20
rect -239 -14 -227 20
rect -285 -48 -227 -14
rect -285 -82 -273 -48
rect -239 -82 -227 -48
rect -285 -116 -227 -82
rect -285 -150 -273 -116
rect -239 -150 -227 -116
rect -285 -184 -227 -150
rect -285 -218 -273 -184
rect -239 -218 -227 -184
rect -285 -252 -227 -218
rect -285 -286 -273 -252
rect -239 -286 -227 -252
rect -285 -320 -227 -286
rect -285 -354 -273 -320
rect -239 -354 -227 -320
rect -285 -381 -227 -354
rect -157 292 -99 319
rect -157 258 -145 292
rect -111 258 -99 292
rect -157 224 -99 258
rect -157 190 -145 224
rect -111 190 -99 224
rect -157 156 -99 190
rect -157 122 -145 156
rect -111 122 -99 156
rect -157 88 -99 122
rect -157 54 -145 88
rect -111 54 -99 88
rect -157 20 -99 54
rect -157 -14 -145 20
rect -111 -14 -99 20
rect -157 -48 -99 -14
rect -157 -82 -145 -48
rect -111 -82 -99 -48
rect -157 -116 -99 -82
rect -157 -150 -145 -116
rect -111 -150 -99 -116
rect -157 -184 -99 -150
rect -157 -218 -145 -184
rect -111 -218 -99 -184
rect -157 -252 -99 -218
rect -157 -286 -145 -252
rect -111 -286 -99 -252
rect -157 -320 -99 -286
rect -157 -354 -145 -320
rect -111 -354 -99 -320
rect -157 -381 -99 -354
rect -29 292 29 319
rect -29 258 -17 292
rect 17 258 29 292
rect -29 224 29 258
rect -29 190 -17 224
rect 17 190 29 224
rect -29 156 29 190
rect -29 122 -17 156
rect 17 122 29 156
rect -29 88 29 122
rect -29 54 -17 88
rect 17 54 29 88
rect -29 20 29 54
rect -29 -14 -17 20
rect 17 -14 29 20
rect -29 -48 29 -14
rect -29 -82 -17 -48
rect 17 -82 29 -48
rect -29 -116 29 -82
rect -29 -150 -17 -116
rect 17 -150 29 -116
rect -29 -184 29 -150
rect -29 -218 -17 -184
rect 17 -218 29 -184
rect -29 -252 29 -218
rect -29 -286 -17 -252
rect 17 -286 29 -252
rect -29 -320 29 -286
rect -29 -354 -17 -320
rect 17 -354 29 -320
rect -29 -381 29 -354
rect 99 292 157 319
rect 99 258 111 292
rect 145 258 157 292
rect 99 224 157 258
rect 99 190 111 224
rect 145 190 157 224
rect 99 156 157 190
rect 99 122 111 156
rect 145 122 157 156
rect 99 88 157 122
rect 99 54 111 88
rect 145 54 157 88
rect 99 20 157 54
rect 99 -14 111 20
rect 145 -14 157 20
rect 99 -48 157 -14
rect 99 -82 111 -48
rect 145 -82 157 -48
rect 99 -116 157 -82
rect 99 -150 111 -116
rect 145 -150 157 -116
rect 99 -184 157 -150
rect 99 -218 111 -184
rect 145 -218 157 -184
rect 99 -252 157 -218
rect 99 -286 111 -252
rect 145 -286 157 -252
rect 99 -320 157 -286
rect 99 -354 111 -320
rect 145 -354 157 -320
rect 99 -381 157 -354
rect 227 292 285 319
rect 227 258 239 292
rect 273 258 285 292
rect 227 224 285 258
rect 227 190 239 224
rect 273 190 285 224
rect 227 156 285 190
rect 227 122 239 156
rect 273 122 285 156
rect 227 88 285 122
rect 227 54 239 88
rect 273 54 285 88
rect 227 20 285 54
rect 227 -14 239 20
rect 273 -14 285 20
rect 227 -48 285 -14
rect 227 -82 239 -48
rect 273 -82 285 -48
rect 227 -116 285 -82
rect 227 -150 239 -116
rect 273 -150 285 -116
rect 227 -184 285 -150
rect 227 -218 239 -184
rect 273 -218 285 -184
rect 227 -252 285 -218
rect 227 -286 239 -252
rect 273 -286 285 -252
rect 227 -320 285 -286
rect 227 -354 239 -320
rect 273 -354 285 -320
rect 227 -381 285 -354
rect 355 292 413 319
rect 355 258 367 292
rect 401 258 413 292
rect 355 224 413 258
rect 355 190 367 224
rect 401 190 413 224
rect 355 156 413 190
rect 355 122 367 156
rect 401 122 413 156
rect 355 88 413 122
rect 355 54 367 88
rect 401 54 413 88
rect 355 20 413 54
rect 355 -14 367 20
rect 401 -14 413 20
rect 355 -48 413 -14
rect 355 -82 367 -48
rect 401 -82 413 -48
rect 355 -116 413 -82
rect 355 -150 367 -116
rect 401 -150 413 -116
rect 355 -184 413 -150
rect 355 -218 367 -184
rect 401 -218 413 -184
rect 355 -252 413 -218
rect 355 -286 367 -252
rect 401 -286 413 -252
rect 355 -320 413 -286
rect 355 -354 367 -320
rect 401 -354 413 -320
rect 355 -381 413 -354
rect 483 292 541 319
rect 483 258 495 292
rect 529 258 541 292
rect 483 224 541 258
rect 483 190 495 224
rect 529 190 541 224
rect 483 156 541 190
rect 483 122 495 156
rect 529 122 541 156
rect 483 88 541 122
rect 483 54 495 88
rect 529 54 541 88
rect 483 20 541 54
rect 483 -14 495 20
rect 529 -14 541 20
rect 483 -48 541 -14
rect 483 -82 495 -48
rect 529 -82 541 -48
rect 483 -116 541 -82
rect 483 -150 495 -116
rect 529 -150 541 -116
rect 483 -184 541 -150
rect 483 -218 495 -184
rect 529 -218 541 -184
rect 483 -252 541 -218
rect 483 -286 495 -252
rect 529 -286 541 -252
rect 483 -320 541 -286
rect 483 -354 495 -320
rect 529 -354 541 -320
rect 483 -381 541 -354
rect 611 292 669 319
rect 611 258 623 292
rect 657 258 669 292
rect 611 224 669 258
rect 611 190 623 224
rect 657 190 669 224
rect 611 156 669 190
rect 611 122 623 156
rect 657 122 669 156
rect 611 88 669 122
rect 611 54 623 88
rect 657 54 669 88
rect 611 20 669 54
rect 611 -14 623 20
rect 657 -14 669 20
rect 611 -48 669 -14
rect 611 -82 623 -48
rect 657 -82 669 -48
rect 611 -116 669 -82
rect 611 -150 623 -116
rect 657 -150 669 -116
rect 611 -184 669 -150
rect 611 -218 623 -184
rect 657 -218 669 -184
rect 611 -252 669 -218
rect 611 -286 623 -252
rect 657 -286 669 -252
rect 611 -320 669 -286
rect 611 -354 623 -320
rect 657 -354 669 -320
rect 611 -381 669 -354
rect 739 292 797 319
rect 739 258 751 292
rect 785 258 797 292
rect 739 224 797 258
rect 739 190 751 224
rect 785 190 797 224
rect 739 156 797 190
rect 739 122 751 156
rect 785 122 797 156
rect 739 88 797 122
rect 739 54 751 88
rect 785 54 797 88
rect 739 20 797 54
rect 739 -14 751 20
rect 785 -14 797 20
rect 739 -48 797 -14
rect 739 -82 751 -48
rect 785 -82 797 -48
rect 739 -116 797 -82
rect 739 -150 751 -116
rect 785 -150 797 -116
rect 739 -184 797 -150
rect 739 -218 751 -184
rect 785 -218 797 -184
rect 739 -252 797 -218
rect 739 -286 751 -252
rect 785 -286 797 -252
rect 739 -320 797 -286
rect 739 -354 751 -320
rect 785 -354 797 -320
rect 739 -381 797 -354
rect 867 292 925 319
rect 867 258 879 292
rect 913 258 925 292
rect 867 224 925 258
rect 867 190 879 224
rect 913 190 925 224
rect 867 156 925 190
rect 867 122 879 156
rect 913 122 925 156
rect 867 88 925 122
rect 867 54 879 88
rect 913 54 925 88
rect 867 20 925 54
rect 867 -14 879 20
rect 913 -14 925 20
rect 867 -48 925 -14
rect 867 -82 879 -48
rect 913 -82 925 -48
rect 867 -116 925 -82
rect 867 -150 879 -116
rect 913 -150 925 -116
rect 867 -184 925 -150
rect 867 -218 879 -184
rect 913 -218 925 -184
rect 867 -252 925 -218
rect 867 -286 879 -252
rect 913 -286 925 -252
rect 867 -320 925 -286
rect 867 -354 879 -320
rect 913 -354 925 -320
rect 867 -381 925 -354
rect 995 292 1053 319
rect 995 258 1007 292
rect 1041 258 1053 292
rect 995 224 1053 258
rect 995 190 1007 224
rect 1041 190 1053 224
rect 995 156 1053 190
rect 995 122 1007 156
rect 1041 122 1053 156
rect 995 88 1053 122
rect 995 54 1007 88
rect 1041 54 1053 88
rect 995 20 1053 54
rect 995 -14 1007 20
rect 1041 -14 1053 20
rect 995 -48 1053 -14
rect 995 -82 1007 -48
rect 1041 -82 1053 -48
rect 995 -116 1053 -82
rect 995 -150 1007 -116
rect 1041 -150 1053 -116
rect 995 -184 1053 -150
rect 995 -218 1007 -184
rect 1041 -218 1053 -184
rect 995 -252 1053 -218
rect 995 -286 1007 -252
rect 1041 -286 1053 -252
rect 995 -320 1053 -286
rect 995 -354 1007 -320
rect 1041 -354 1053 -320
rect 995 -381 1053 -354
rect 1123 292 1181 319
rect 1123 258 1135 292
rect 1169 258 1181 292
rect 1123 224 1181 258
rect 1123 190 1135 224
rect 1169 190 1181 224
rect 1123 156 1181 190
rect 1123 122 1135 156
rect 1169 122 1181 156
rect 1123 88 1181 122
rect 1123 54 1135 88
rect 1169 54 1181 88
rect 1123 20 1181 54
rect 1123 -14 1135 20
rect 1169 -14 1181 20
rect 1123 -48 1181 -14
rect 1123 -82 1135 -48
rect 1169 -82 1181 -48
rect 1123 -116 1181 -82
rect 1123 -150 1135 -116
rect 1169 -150 1181 -116
rect 1123 -184 1181 -150
rect 1123 -218 1135 -184
rect 1169 -218 1181 -184
rect 1123 -252 1181 -218
rect 1123 -286 1135 -252
rect 1169 -286 1181 -252
rect 1123 -320 1181 -286
rect 1123 -354 1135 -320
rect 1169 -354 1181 -320
rect 1123 -381 1181 -354
rect 1251 292 1309 319
rect 1251 258 1263 292
rect 1297 258 1309 292
rect 1251 224 1309 258
rect 1251 190 1263 224
rect 1297 190 1309 224
rect 1251 156 1309 190
rect 1251 122 1263 156
rect 1297 122 1309 156
rect 1251 88 1309 122
rect 1251 54 1263 88
rect 1297 54 1309 88
rect 1251 20 1309 54
rect 1251 -14 1263 20
rect 1297 -14 1309 20
rect 1251 -48 1309 -14
rect 1251 -82 1263 -48
rect 1297 -82 1309 -48
rect 1251 -116 1309 -82
rect 1251 -150 1263 -116
rect 1297 -150 1309 -116
rect 1251 -184 1309 -150
rect 1251 -218 1263 -184
rect 1297 -218 1309 -184
rect 1251 -252 1309 -218
rect 1251 -286 1263 -252
rect 1297 -286 1309 -252
rect 1251 -320 1309 -286
rect 1251 -354 1263 -320
rect 1297 -354 1309 -320
rect 1251 -381 1309 -354
rect 1379 292 1437 319
rect 1379 258 1391 292
rect 1425 258 1437 292
rect 1379 224 1437 258
rect 1379 190 1391 224
rect 1425 190 1437 224
rect 1379 156 1437 190
rect 1379 122 1391 156
rect 1425 122 1437 156
rect 1379 88 1437 122
rect 1379 54 1391 88
rect 1425 54 1437 88
rect 1379 20 1437 54
rect 1379 -14 1391 20
rect 1425 -14 1437 20
rect 1379 -48 1437 -14
rect 1379 -82 1391 -48
rect 1425 -82 1437 -48
rect 1379 -116 1437 -82
rect 1379 -150 1391 -116
rect 1425 -150 1437 -116
rect 1379 -184 1437 -150
rect 1379 -218 1391 -184
rect 1425 -218 1437 -184
rect 1379 -252 1437 -218
rect 1379 -286 1391 -252
rect 1425 -286 1437 -252
rect 1379 -320 1437 -286
rect 1379 -354 1391 -320
rect 1425 -354 1437 -320
rect 1379 -381 1437 -354
rect 1507 292 1565 319
rect 1507 258 1519 292
rect 1553 258 1565 292
rect 1507 224 1565 258
rect 1507 190 1519 224
rect 1553 190 1565 224
rect 1507 156 1565 190
rect 1507 122 1519 156
rect 1553 122 1565 156
rect 1507 88 1565 122
rect 1507 54 1519 88
rect 1553 54 1565 88
rect 1507 20 1565 54
rect 1507 -14 1519 20
rect 1553 -14 1565 20
rect 1507 -48 1565 -14
rect 1507 -82 1519 -48
rect 1553 -82 1565 -48
rect 1507 -116 1565 -82
rect 1507 -150 1519 -116
rect 1553 -150 1565 -116
rect 1507 -184 1565 -150
rect 1507 -218 1519 -184
rect 1553 -218 1565 -184
rect 1507 -252 1565 -218
rect 1507 -286 1519 -252
rect 1553 -286 1565 -252
rect 1507 -320 1565 -286
rect 1507 -354 1519 -320
rect 1553 -354 1565 -320
rect 1507 -381 1565 -354
rect 1635 292 1693 319
rect 1635 258 1647 292
rect 1681 258 1693 292
rect 1635 224 1693 258
rect 1635 190 1647 224
rect 1681 190 1693 224
rect 1635 156 1693 190
rect 1635 122 1647 156
rect 1681 122 1693 156
rect 1635 88 1693 122
rect 1635 54 1647 88
rect 1681 54 1693 88
rect 1635 20 1693 54
rect 1635 -14 1647 20
rect 1681 -14 1693 20
rect 1635 -48 1693 -14
rect 1635 -82 1647 -48
rect 1681 -82 1693 -48
rect 1635 -116 1693 -82
rect 1635 -150 1647 -116
rect 1681 -150 1693 -116
rect 1635 -184 1693 -150
rect 1635 -218 1647 -184
rect 1681 -218 1693 -184
rect 1635 -252 1693 -218
rect 1635 -286 1647 -252
rect 1681 -286 1693 -252
rect 1635 -320 1693 -286
rect 1635 -354 1647 -320
rect 1681 -354 1693 -320
rect 1635 -381 1693 -354
rect 1763 292 1821 319
rect 1763 258 1775 292
rect 1809 258 1821 292
rect 1763 224 1821 258
rect 1763 190 1775 224
rect 1809 190 1821 224
rect 1763 156 1821 190
rect 1763 122 1775 156
rect 1809 122 1821 156
rect 1763 88 1821 122
rect 1763 54 1775 88
rect 1809 54 1821 88
rect 1763 20 1821 54
rect 1763 -14 1775 20
rect 1809 -14 1821 20
rect 1763 -48 1821 -14
rect 1763 -82 1775 -48
rect 1809 -82 1821 -48
rect 1763 -116 1821 -82
rect 1763 -150 1775 -116
rect 1809 -150 1821 -116
rect 1763 -184 1821 -150
rect 1763 -218 1775 -184
rect 1809 -218 1821 -184
rect 1763 -252 1821 -218
rect 1763 -286 1775 -252
rect 1809 -286 1821 -252
rect 1763 -320 1821 -286
rect 1763 -354 1775 -320
rect 1809 -354 1821 -320
rect 1763 -381 1821 -354
rect 1891 292 1949 319
rect 1891 258 1903 292
rect 1937 258 1949 292
rect 1891 224 1949 258
rect 1891 190 1903 224
rect 1937 190 1949 224
rect 1891 156 1949 190
rect 1891 122 1903 156
rect 1937 122 1949 156
rect 1891 88 1949 122
rect 1891 54 1903 88
rect 1937 54 1949 88
rect 1891 20 1949 54
rect 1891 -14 1903 20
rect 1937 -14 1949 20
rect 1891 -48 1949 -14
rect 1891 -82 1903 -48
rect 1937 -82 1949 -48
rect 1891 -116 1949 -82
rect 1891 -150 1903 -116
rect 1937 -150 1949 -116
rect 1891 -184 1949 -150
rect 1891 -218 1903 -184
rect 1937 -218 1949 -184
rect 1891 -252 1949 -218
rect 1891 -286 1903 -252
rect 1937 -286 1949 -252
rect 1891 -320 1949 -286
rect 1891 -354 1903 -320
rect 1937 -354 1949 -320
rect 1891 -381 1949 -354
rect 2019 292 2077 319
rect 2019 258 2031 292
rect 2065 258 2077 292
rect 2019 224 2077 258
rect 2019 190 2031 224
rect 2065 190 2077 224
rect 2019 156 2077 190
rect 2019 122 2031 156
rect 2065 122 2077 156
rect 2019 88 2077 122
rect 2019 54 2031 88
rect 2065 54 2077 88
rect 2019 20 2077 54
rect 2019 -14 2031 20
rect 2065 -14 2077 20
rect 2019 -48 2077 -14
rect 2019 -82 2031 -48
rect 2065 -82 2077 -48
rect 2019 -116 2077 -82
rect 2019 -150 2031 -116
rect 2065 -150 2077 -116
rect 2019 -184 2077 -150
rect 2019 -218 2031 -184
rect 2065 -218 2077 -184
rect 2019 -252 2077 -218
rect 2019 -286 2031 -252
rect 2065 -286 2077 -252
rect 2019 -320 2077 -286
rect 2019 -354 2031 -320
rect 2065 -354 2077 -320
rect 2019 -381 2077 -354
<< ndiffc >>
rect -2065 258 -2031 292
rect -2065 190 -2031 224
rect -2065 122 -2031 156
rect -2065 54 -2031 88
rect -2065 -14 -2031 20
rect -2065 -82 -2031 -48
rect -2065 -150 -2031 -116
rect -2065 -218 -2031 -184
rect -2065 -286 -2031 -252
rect -2065 -354 -2031 -320
rect -1937 258 -1903 292
rect -1937 190 -1903 224
rect -1937 122 -1903 156
rect -1937 54 -1903 88
rect -1937 -14 -1903 20
rect -1937 -82 -1903 -48
rect -1937 -150 -1903 -116
rect -1937 -218 -1903 -184
rect -1937 -286 -1903 -252
rect -1937 -354 -1903 -320
rect -1809 258 -1775 292
rect -1809 190 -1775 224
rect -1809 122 -1775 156
rect -1809 54 -1775 88
rect -1809 -14 -1775 20
rect -1809 -82 -1775 -48
rect -1809 -150 -1775 -116
rect -1809 -218 -1775 -184
rect -1809 -286 -1775 -252
rect -1809 -354 -1775 -320
rect -1681 258 -1647 292
rect -1681 190 -1647 224
rect -1681 122 -1647 156
rect -1681 54 -1647 88
rect -1681 -14 -1647 20
rect -1681 -82 -1647 -48
rect -1681 -150 -1647 -116
rect -1681 -218 -1647 -184
rect -1681 -286 -1647 -252
rect -1681 -354 -1647 -320
rect -1553 258 -1519 292
rect -1553 190 -1519 224
rect -1553 122 -1519 156
rect -1553 54 -1519 88
rect -1553 -14 -1519 20
rect -1553 -82 -1519 -48
rect -1553 -150 -1519 -116
rect -1553 -218 -1519 -184
rect -1553 -286 -1519 -252
rect -1553 -354 -1519 -320
rect -1425 258 -1391 292
rect -1425 190 -1391 224
rect -1425 122 -1391 156
rect -1425 54 -1391 88
rect -1425 -14 -1391 20
rect -1425 -82 -1391 -48
rect -1425 -150 -1391 -116
rect -1425 -218 -1391 -184
rect -1425 -286 -1391 -252
rect -1425 -354 -1391 -320
rect -1297 258 -1263 292
rect -1297 190 -1263 224
rect -1297 122 -1263 156
rect -1297 54 -1263 88
rect -1297 -14 -1263 20
rect -1297 -82 -1263 -48
rect -1297 -150 -1263 -116
rect -1297 -218 -1263 -184
rect -1297 -286 -1263 -252
rect -1297 -354 -1263 -320
rect -1169 258 -1135 292
rect -1169 190 -1135 224
rect -1169 122 -1135 156
rect -1169 54 -1135 88
rect -1169 -14 -1135 20
rect -1169 -82 -1135 -48
rect -1169 -150 -1135 -116
rect -1169 -218 -1135 -184
rect -1169 -286 -1135 -252
rect -1169 -354 -1135 -320
rect -1041 258 -1007 292
rect -1041 190 -1007 224
rect -1041 122 -1007 156
rect -1041 54 -1007 88
rect -1041 -14 -1007 20
rect -1041 -82 -1007 -48
rect -1041 -150 -1007 -116
rect -1041 -218 -1007 -184
rect -1041 -286 -1007 -252
rect -1041 -354 -1007 -320
rect -913 258 -879 292
rect -913 190 -879 224
rect -913 122 -879 156
rect -913 54 -879 88
rect -913 -14 -879 20
rect -913 -82 -879 -48
rect -913 -150 -879 -116
rect -913 -218 -879 -184
rect -913 -286 -879 -252
rect -913 -354 -879 -320
rect -785 258 -751 292
rect -785 190 -751 224
rect -785 122 -751 156
rect -785 54 -751 88
rect -785 -14 -751 20
rect -785 -82 -751 -48
rect -785 -150 -751 -116
rect -785 -218 -751 -184
rect -785 -286 -751 -252
rect -785 -354 -751 -320
rect -657 258 -623 292
rect -657 190 -623 224
rect -657 122 -623 156
rect -657 54 -623 88
rect -657 -14 -623 20
rect -657 -82 -623 -48
rect -657 -150 -623 -116
rect -657 -218 -623 -184
rect -657 -286 -623 -252
rect -657 -354 -623 -320
rect -529 258 -495 292
rect -529 190 -495 224
rect -529 122 -495 156
rect -529 54 -495 88
rect -529 -14 -495 20
rect -529 -82 -495 -48
rect -529 -150 -495 -116
rect -529 -218 -495 -184
rect -529 -286 -495 -252
rect -529 -354 -495 -320
rect -401 258 -367 292
rect -401 190 -367 224
rect -401 122 -367 156
rect -401 54 -367 88
rect -401 -14 -367 20
rect -401 -82 -367 -48
rect -401 -150 -367 -116
rect -401 -218 -367 -184
rect -401 -286 -367 -252
rect -401 -354 -367 -320
rect -273 258 -239 292
rect -273 190 -239 224
rect -273 122 -239 156
rect -273 54 -239 88
rect -273 -14 -239 20
rect -273 -82 -239 -48
rect -273 -150 -239 -116
rect -273 -218 -239 -184
rect -273 -286 -239 -252
rect -273 -354 -239 -320
rect -145 258 -111 292
rect -145 190 -111 224
rect -145 122 -111 156
rect -145 54 -111 88
rect -145 -14 -111 20
rect -145 -82 -111 -48
rect -145 -150 -111 -116
rect -145 -218 -111 -184
rect -145 -286 -111 -252
rect -145 -354 -111 -320
rect -17 258 17 292
rect -17 190 17 224
rect -17 122 17 156
rect -17 54 17 88
rect -17 -14 17 20
rect -17 -82 17 -48
rect -17 -150 17 -116
rect -17 -218 17 -184
rect -17 -286 17 -252
rect -17 -354 17 -320
rect 111 258 145 292
rect 111 190 145 224
rect 111 122 145 156
rect 111 54 145 88
rect 111 -14 145 20
rect 111 -82 145 -48
rect 111 -150 145 -116
rect 111 -218 145 -184
rect 111 -286 145 -252
rect 111 -354 145 -320
rect 239 258 273 292
rect 239 190 273 224
rect 239 122 273 156
rect 239 54 273 88
rect 239 -14 273 20
rect 239 -82 273 -48
rect 239 -150 273 -116
rect 239 -218 273 -184
rect 239 -286 273 -252
rect 239 -354 273 -320
rect 367 258 401 292
rect 367 190 401 224
rect 367 122 401 156
rect 367 54 401 88
rect 367 -14 401 20
rect 367 -82 401 -48
rect 367 -150 401 -116
rect 367 -218 401 -184
rect 367 -286 401 -252
rect 367 -354 401 -320
rect 495 258 529 292
rect 495 190 529 224
rect 495 122 529 156
rect 495 54 529 88
rect 495 -14 529 20
rect 495 -82 529 -48
rect 495 -150 529 -116
rect 495 -218 529 -184
rect 495 -286 529 -252
rect 495 -354 529 -320
rect 623 258 657 292
rect 623 190 657 224
rect 623 122 657 156
rect 623 54 657 88
rect 623 -14 657 20
rect 623 -82 657 -48
rect 623 -150 657 -116
rect 623 -218 657 -184
rect 623 -286 657 -252
rect 623 -354 657 -320
rect 751 258 785 292
rect 751 190 785 224
rect 751 122 785 156
rect 751 54 785 88
rect 751 -14 785 20
rect 751 -82 785 -48
rect 751 -150 785 -116
rect 751 -218 785 -184
rect 751 -286 785 -252
rect 751 -354 785 -320
rect 879 258 913 292
rect 879 190 913 224
rect 879 122 913 156
rect 879 54 913 88
rect 879 -14 913 20
rect 879 -82 913 -48
rect 879 -150 913 -116
rect 879 -218 913 -184
rect 879 -286 913 -252
rect 879 -354 913 -320
rect 1007 258 1041 292
rect 1007 190 1041 224
rect 1007 122 1041 156
rect 1007 54 1041 88
rect 1007 -14 1041 20
rect 1007 -82 1041 -48
rect 1007 -150 1041 -116
rect 1007 -218 1041 -184
rect 1007 -286 1041 -252
rect 1007 -354 1041 -320
rect 1135 258 1169 292
rect 1135 190 1169 224
rect 1135 122 1169 156
rect 1135 54 1169 88
rect 1135 -14 1169 20
rect 1135 -82 1169 -48
rect 1135 -150 1169 -116
rect 1135 -218 1169 -184
rect 1135 -286 1169 -252
rect 1135 -354 1169 -320
rect 1263 258 1297 292
rect 1263 190 1297 224
rect 1263 122 1297 156
rect 1263 54 1297 88
rect 1263 -14 1297 20
rect 1263 -82 1297 -48
rect 1263 -150 1297 -116
rect 1263 -218 1297 -184
rect 1263 -286 1297 -252
rect 1263 -354 1297 -320
rect 1391 258 1425 292
rect 1391 190 1425 224
rect 1391 122 1425 156
rect 1391 54 1425 88
rect 1391 -14 1425 20
rect 1391 -82 1425 -48
rect 1391 -150 1425 -116
rect 1391 -218 1425 -184
rect 1391 -286 1425 -252
rect 1391 -354 1425 -320
rect 1519 258 1553 292
rect 1519 190 1553 224
rect 1519 122 1553 156
rect 1519 54 1553 88
rect 1519 -14 1553 20
rect 1519 -82 1553 -48
rect 1519 -150 1553 -116
rect 1519 -218 1553 -184
rect 1519 -286 1553 -252
rect 1519 -354 1553 -320
rect 1647 258 1681 292
rect 1647 190 1681 224
rect 1647 122 1681 156
rect 1647 54 1681 88
rect 1647 -14 1681 20
rect 1647 -82 1681 -48
rect 1647 -150 1681 -116
rect 1647 -218 1681 -184
rect 1647 -286 1681 -252
rect 1647 -354 1681 -320
rect 1775 258 1809 292
rect 1775 190 1809 224
rect 1775 122 1809 156
rect 1775 54 1809 88
rect 1775 -14 1809 20
rect 1775 -82 1809 -48
rect 1775 -150 1809 -116
rect 1775 -218 1809 -184
rect 1775 -286 1809 -252
rect 1775 -354 1809 -320
rect 1903 258 1937 292
rect 1903 190 1937 224
rect 1903 122 1937 156
rect 1903 54 1937 88
rect 1903 -14 1937 20
rect 1903 -82 1937 -48
rect 1903 -150 1937 -116
rect 1903 -218 1937 -184
rect 1903 -286 1937 -252
rect 1903 -354 1937 -320
rect 2031 258 2065 292
rect 2031 190 2065 224
rect 2031 122 2065 156
rect 2031 54 2065 88
rect 2031 -14 2065 20
rect 2031 -82 2065 -48
rect 2031 -150 2065 -116
rect 2031 -218 2065 -184
rect 2031 -286 2065 -252
rect 2031 -354 2065 -320
<< psubdiff >>
rect -2179 459 -2057 493
rect -2023 459 -1989 493
rect -1955 459 -1921 493
rect -1887 459 -1853 493
rect -1819 459 -1785 493
rect -1751 459 -1717 493
rect -1683 459 -1649 493
rect -1615 459 -1581 493
rect -1547 459 -1513 493
rect -1479 459 -1445 493
rect -1411 459 -1377 493
rect -1343 459 -1309 493
rect -1275 459 -1241 493
rect -1207 459 -1173 493
rect -1139 459 -1105 493
rect -1071 459 -1037 493
rect -1003 459 -969 493
rect -935 459 -901 493
rect -867 459 -833 493
rect -799 459 -765 493
rect -731 459 -697 493
rect -663 459 -629 493
rect -595 459 -561 493
rect -527 459 -493 493
rect -459 459 -425 493
rect -391 459 -357 493
rect -323 459 -289 493
rect -255 459 -221 493
rect -187 459 -153 493
rect -119 459 -85 493
rect -51 459 -17 493
rect 17 459 51 493
rect 85 459 119 493
rect 153 459 187 493
rect 221 459 255 493
rect 289 459 323 493
rect 357 459 391 493
rect 425 459 459 493
rect 493 459 527 493
rect 561 459 595 493
rect 629 459 663 493
rect 697 459 731 493
rect 765 459 799 493
rect 833 459 867 493
rect 901 459 935 493
rect 969 459 1003 493
rect 1037 459 1071 493
rect 1105 459 1139 493
rect 1173 459 1207 493
rect 1241 459 1275 493
rect 1309 459 1343 493
rect 1377 459 1411 493
rect 1445 459 1479 493
rect 1513 459 1547 493
rect 1581 459 1615 493
rect 1649 459 1683 493
rect 1717 459 1751 493
rect 1785 459 1819 493
rect 1853 459 1887 493
rect 1921 459 1955 493
rect 1989 459 2023 493
rect 2057 459 2179 493
rect -2179 391 -2145 459
rect -2179 323 -2145 357
rect 2145 391 2179 459
rect 2145 323 2179 357
rect -2179 255 -2145 289
rect -2179 187 -2145 221
rect -2179 119 -2145 153
rect -2179 51 -2145 85
rect -2179 -17 -2145 17
rect -2179 -85 -2145 -51
rect -2179 -153 -2145 -119
rect -2179 -221 -2145 -187
rect -2179 -289 -2145 -255
rect -2179 -357 -2145 -323
rect 2145 255 2179 289
rect 2145 187 2179 221
rect 2145 119 2179 153
rect 2145 51 2179 85
rect 2145 -17 2179 17
rect 2145 -85 2179 -51
rect 2145 -153 2179 -119
rect 2145 -221 2179 -187
rect 2145 -289 2179 -255
rect 2145 -357 2179 -323
rect -2179 -459 -2145 -391
rect 2145 -459 2179 -391
rect -2179 -493 -2057 -459
rect -2023 -493 -1989 -459
rect -1955 -493 -1921 -459
rect -1887 -493 -1853 -459
rect -1819 -493 -1785 -459
rect -1751 -493 -1717 -459
rect -1683 -493 -1649 -459
rect -1615 -493 -1581 -459
rect -1547 -493 -1513 -459
rect -1479 -493 -1445 -459
rect -1411 -493 -1377 -459
rect -1343 -493 -1309 -459
rect -1275 -493 -1241 -459
rect -1207 -493 -1173 -459
rect -1139 -493 -1105 -459
rect -1071 -493 -1037 -459
rect -1003 -493 -969 -459
rect -935 -493 -901 -459
rect -867 -493 -833 -459
rect -799 -493 -765 -459
rect -731 -493 -697 -459
rect -663 -493 -629 -459
rect -595 -493 -561 -459
rect -527 -493 -493 -459
rect -459 -493 -425 -459
rect -391 -493 -357 -459
rect -323 -493 -289 -459
rect -255 -493 -221 -459
rect -187 -493 -153 -459
rect -119 -493 -85 -459
rect -51 -493 -17 -459
rect 17 -493 51 -459
rect 85 -493 119 -459
rect 153 -493 187 -459
rect 221 -493 255 -459
rect 289 -493 323 -459
rect 357 -493 391 -459
rect 425 -493 459 -459
rect 493 -493 527 -459
rect 561 -493 595 -459
rect 629 -493 663 -459
rect 697 -493 731 -459
rect 765 -493 799 -459
rect 833 -493 867 -459
rect 901 -493 935 -459
rect 969 -493 1003 -459
rect 1037 -493 1071 -459
rect 1105 -493 1139 -459
rect 1173 -493 1207 -459
rect 1241 -493 1275 -459
rect 1309 -493 1343 -459
rect 1377 -493 1411 -459
rect 1445 -493 1479 -459
rect 1513 -493 1547 -459
rect 1581 -493 1615 -459
rect 1649 -493 1683 -459
rect 1717 -493 1751 -459
rect 1785 -493 1819 -459
rect 1853 -493 1887 -459
rect 1921 -493 1955 -459
rect 1989 -493 2023 -459
rect 2057 -493 2179 -459
<< psubdiffcont >>
rect -2057 459 -2023 493
rect -1989 459 -1955 493
rect -1921 459 -1887 493
rect -1853 459 -1819 493
rect -1785 459 -1751 493
rect -1717 459 -1683 493
rect -1649 459 -1615 493
rect -1581 459 -1547 493
rect -1513 459 -1479 493
rect -1445 459 -1411 493
rect -1377 459 -1343 493
rect -1309 459 -1275 493
rect -1241 459 -1207 493
rect -1173 459 -1139 493
rect -1105 459 -1071 493
rect -1037 459 -1003 493
rect -969 459 -935 493
rect -901 459 -867 493
rect -833 459 -799 493
rect -765 459 -731 493
rect -697 459 -663 493
rect -629 459 -595 493
rect -561 459 -527 493
rect -493 459 -459 493
rect -425 459 -391 493
rect -357 459 -323 493
rect -289 459 -255 493
rect -221 459 -187 493
rect -153 459 -119 493
rect -85 459 -51 493
rect -17 459 17 493
rect 51 459 85 493
rect 119 459 153 493
rect 187 459 221 493
rect 255 459 289 493
rect 323 459 357 493
rect 391 459 425 493
rect 459 459 493 493
rect 527 459 561 493
rect 595 459 629 493
rect 663 459 697 493
rect 731 459 765 493
rect 799 459 833 493
rect 867 459 901 493
rect 935 459 969 493
rect 1003 459 1037 493
rect 1071 459 1105 493
rect 1139 459 1173 493
rect 1207 459 1241 493
rect 1275 459 1309 493
rect 1343 459 1377 493
rect 1411 459 1445 493
rect 1479 459 1513 493
rect 1547 459 1581 493
rect 1615 459 1649 493
rect 1683 459 1717 493
rect 1751 459 1785 493
rect 1819 459 1853 493
rect 1887 459 1921 493
rect 1955 459 1989 493
rect 2023 459 2057 493
rect -2179 357 -2145 391
rect -2179 289 -2145 323
rect 2145 357 2179 391
rect -2179 221 -2145 255
rect -2179 153 -2145 187
rect -2179 85 -2145 119
rect -2179 17 -2145 51
rect -2179 -51 -2145 -17
rect -2179 -119 -2145 -85
rect -2179 -187 -2145 -153
rect -2179 -255 -2145 -221
rect -2179 -323 -2145 -289
rect -2179 -391 -2145 -357
rect 2145 289 2179 323
rect 2145 221 2179 255
rect 2145 153 2179 187
rect 2145 85 2179 119
rect 2145 17 2179 51
rect 2145 -51 2179 -17
rect 2145 -119 2179 -85
rect 2145 -187 2179 -153
rect 2145 -255 2179 -221
rect 2145 -323 2179 -289
rect 2145 -391 2179 -357
rect -2057 -493 -2023 -459
rect -1989 -493 -1955 -459
rect -1921 -493 -1887 -459
rect -1853 -493 -1819 -459
rect -1785 -493 -1751 -459
rect -1717 -493 -1683 -459
rect -1649 -493 -1615 -459
rect -1581 -493 -1547 -459
rect -1513 -493 -1479 -459
rect -1445 -493 -1411 -459
rect -1377 -493 -1343 -459
rect -1309 -493 -1275 -459
rect -1241 -493 -1207 -459
rect -1173 -493 -1139 -459
rect -1105 -493 -1071 -459
rect -1037 -493 -1003 -459
rect -969 -493 -935 -459
rect -901 -493 -867 -459
rect -833 -493 -799 -459
rect -765 -493 -731 -459
rect -697 -493 -663 -459
rect -629 -493 -595 -459
rect -561 -493 -527 -459
rect -493 -493 -459 -459
rect -425 -493 -391 -459
rect -357 -493 -323 -459
rect -289 -493 -255 -459
rect -221 -493 -187 -459
rect -153 -493 -119 -459
rect -85 -493 -51 -459
rect -17 -493 17 -459
rect 51 -493 85 -459
rect 119 -493 153 -459
rect 187 -493 221 -459
rect 255 -493 289 -459
rect 323 -493 357 -459
rect 391 -493 425 -459
rect 459 -493 493 -459
rect 527 -493 561 -459
rect 595 -493 629 -459
rect 663 -493 697 -459
rect 731 -493 765 -459
rect 799 -493 833 -459
rect 867 -493 901 -459
rect 935 -493 969 -459
rect 1003 -493 1037 -459
rect 1071 -493 1105 -459
rect 1139 -493 1173 -459
rect 1207 -493 1241 -459
rect 1275 -493 1309 -459
rect 1343 -493 1377 -459
rect 1411 -493 1445 -459
rect 1479 -493 1513 -459
rect 1547 -493 1581 -459
rect 1615 -493 1649 -459
rect 1683 -493 1717 -459
rect 1751 -493 1785 -459
rect 1819 -493 1853 -459
rect 1887 -493 1921 -459
rect 1955 -493 1989 -459
rect 2023 -493 2057 -459
<< poly >>
rect -2019 391 -1949 407
rect -2019 357 -2001 391
rect -1967 357 -1949 391
rect -2019 319 -1949 357
rect -1891 391 -1821 407
rect -1891 357 -1873 391
rect -1839 357 -1821 391
rect -1891 319 -1821 357
rect -1763 391 -1693 407
rect -1763 357 -1745 391
rect -1711 357 -1693 391
rect -1763 319 -1693 357
rect -1635 391 -1565 407
rect -1635 357 -1617 391
rect -1583 357 -1565 391
rect -1635 319 -1565 357
rect -1507 391 -1437 407
rect -1507 357 -1489 391
rect -1455 357 -1437 391
rect -1507 319 -1437 357
rect -1379 391 -1309 407
rect -1379 357 -1361 391
rect -1327 357 -1309 391
rect -1379 319 -1309 357
rect -1251 391 -1181 407
rect -1251 357 -1233 391
rect -1199 357 -1181 391
rect -1251 319 -1181 357
rect -1123 391 -1053 407
rect -1123 357 -1105 391
rect -1071 357 -1053 391
rect -1123 319 -1053 357
rect -995 391 -925 407
rect -995 357 -977 391
rect -943 357 -925 391
rect -995 319 -925 357
rect -867 391 -797 407
rect -867 357 -849 391
rect -815 357 -797 391
rect -867 319 -797 357
rect -739 391 -669 407
rect -739 357 -721 391
rect -687 357 -669 391
rect -739 319 -669 357
rect -611 391 -541 407
rect -611 357 -593 391
rect -559 357 -541 391
rect -611 319 -541 357
rect -483 391 -413 407
rect -483 357 -465 391
rect -431 357 -413 391
rect -483 319 -413 357
rect -355 391 -285 407
rect -355 357 -337 391
rect -303 357 -285 391
rect -355 319 -285 357
rect -227 391 -157 407
rect -227 357 -209 391
rect -175 357 -157 391
rect -227 319 -157 357
rect -99 391 -29 407
rect -99 357 -81 391
rect -47 357 -29 391
rect -99 319 -29 357
rect 29 391 99 407
rect 29 357 47 391
rect 81 357 99 391
rect 29 319 99 357
rect 157 391 227 407
rect 157 357 175 391
rect 209 357 227 391
rect 157 319 227 357
rect 285 391 355 407
rect 285 357 303 391
rect 337 357 355 391
rect 285 319 355 357
rect 413 391 483 407
rect 413 357 431 391
rect 465 357 483 391
rect 413 319 483 357
rect 541 391 611 407
rect 541 357 559 391
rect 593 357 611 391
rect 541 319 611 357
rect 669 391 739 407
rect 669 357 687 391
rect 721 357 739 391
rect 669 319 739 357
rect 797 391 867 407
rect 797 357 815 391
rect 849 357 867 391
rect 797 319 867 357
rect 925 391 995 407
rect 925 357 943 391
rect 977 357 995 391
rect 925 319 995 357
rect 1053 391 1123 407
rect 1053 357 1071 391
rect 1105 357 1123 391
rect 1053 319 1123 357
rect 1181 391 1251 407
rect 1181 357 1199 391
rect 1233 357 1251 391
rect 1181 319 1251 357
rect 1309 391 1379 407
rect 1309 357 1327 391
rect 1361 357 1379 391
rect 1309 319 1379 357
rect 1437 391 1507 407
rect 1437 357 1455 391
rect 1489 357 1507 391
rect 1437 319 1507 357
rect 1565 391 1635 407
rect 1565 357 1583 391
rect 1617 357 1635 391
rect 1565 319 1635 357
rect 1693 391 1763 407
rect 1693 357 1711 391
rect 1745 357 1763 391
rect 1693 319 1763 357
rect 1821 391 1891 407
rect 1821 357 1839 391
rect 1873 357 1891 391
rect 1821 319 1891 357
rect 1949 391 2019 407
rect 1949 357 1967 391
rect 2001 357 2019 391
rect 1949 319 2019 357
rect -2019 -407 -1949 -381
rect -1891 -407 -1821 -381
rect -1763 -407 -1693 -381
rect -1635 -407 -1565 -381
rect -1507 -407 -1437 -381
rect -1379 -407 -1309 -381
rect -1251 -407 -1181 -381
rect -1123 -407 -1053 -381
rect -995 -407 -925 -381
rect -867 -407 -797 -381
rect -739 -407 -669 -381
rect -611 -407 -541 -381
rect -483 -407 -413 -381
rect -355 -407 -285 -381
rect -227 -407 -157 -381
rect -99 -407 -29 -381
rect 29 -407 99 -381
rect 157 -407 227 -381
rect 285 -407 355 -381
rect 413 -407 483 -381
rect 541 -407 611 -381
rect 669 -407 739 -381
rect 797 -407 867 -381
rect 925 -407 995 -381
rect 1053 -407 1123 -381
rect 1181 -407 1251 -381
rect 1309 -407 1379 -381
rect 1437 -407 1507 -381
rect 1565 -407 1635 -381
rect 1693 -407 1763 -381
rect 1821 -407 1891 -381
rect 1949 -407 2019 -381
<< polycont >>
rect -2001 357 -1967 391
rect -1873 357 -1839 391
rect -1745 357 -1711 391
rect -1617 357 -1583 391
rect -1489 357 -1455 391
rect -1361 357 -1327 391
rect -1233 357 -1199 391
rect -1105 357 -1071 391
rect -977 357 -943 391
rect -849 357 -815 391
rect -721 357 -687 391
rect -593 357 -559 391
rect -465 357 -431 391
rect -337 357 -303 391
rect -209 357 -175 391
rect -81 357 -47 391
rect 47 357 81 391
rect 175 357 209 391
rect 303 357 337 391
rect 431 357 465 391
rect 559 357 593 391
rect 687 357 721 391
rect 815 357 849 391
rect 943 357 977 391
rect 1071 357 1105 391
rect 1199 357 1233 391
rect 1327 357 1361 391
rect 1455 357 1489 391
rect 1583 357 1617 391
rect 1711 357 1745 391
rect 1839 357 1873 391
rect 1967 357 2001 391
<< locali >>
rect -2179 459 -2057 493
rect -2023 459 -1989 493
rect -1955 459 -1921 493
rect -1887 459 -1853 493
rect -1819 459 -1785 493
rect -1751 459 -1717 493
rect -1683 459 -1649 493
rect -1615 459 -1581 493
rect -1547 459 -1513 493
rect -1479 459 -1445 493
rect -1411 459 -1377 493
rect -1343 459 -1309 493
rect -1275 459 -1241 493
rect -1207 459 -1173 493
rect -1139 459 -1105 493
rect -1071 459 -1037 493
rect -1003 459 -969 493
rect -935 459 -901 493
rect -867 459 -833 493
rect -799 459 -765 493
rect -731 459 -697 493
rect -663 459 -629 493
rect -595 459 -561 493
rect -527 459 -493 493
rect -459 459 -425 493
rect -391 459 -357 493
rect -323 459 -289 493
rect -255 459 -221 493
rect -187 459 -153 493
rect -119 459 -85 493
rect -51 459 -17 493
rect 17 459 51 493
rect 85 459 119 493
rect 153 459 187 493
rect 221 459 255 493
rect 289 459 323 493
rect 357 459 391 493
rect 425 459 459 493
rect 493 459 527 493
rect 561 459 595 493
rect 629 459 663 493
rect 697 459 731 493
rect 765 459 799 493
rect 833 459 867 493
rect 901 459 935 493
rect 969 459 1003 493
rect 1037 459 1071 493
rect 1105 459 1139 493
rect 1173 459 1207 493
rect 1241 459 1275 493
rect 1309 459 1343 493
rect 1377 459 1411 493
rect 1445 459 1479 493
rect 1513 459 1547 493
rect 1581 459 1615 493
rect 1649 459 1683 493
rect 1717 459 1751 493
rect 1785 459 1819 493
rect 1853 459 1887 493
rect 1921 459 1955 493
rect 1989 459 2023 493
rect 2057 459 2179 493
rect -2179 391 -2145 459
rect 2145 391 2179 459
rect -2019 357 -2001 391
rect -1967 357 -1949 391
rect -1891 357 -1873 391
rect -1839 357 -1821 391
rect -1763 357 -1745 391
rect -1711 357 -1693 391
rect -1635 357 -1617 391
rect -1583 357 -1565 391
rect -1507 357 -1489 391
rect -1455 357 -1437 391
rect -1379 357 -1361 391
rect -1327 357 -1309 391
rect -1251 357 -1233 391
rect -1199 357 -1181 391
rect -1123 357 -1105 391
rect -1071 357 -1053 391
rect -995 357 -977 391
rect -943 357 -925 391
rect -867 357 -849 391
rect -815 357 -797 391
rect -739 357 -721 391
rect -687 357 -669 391
rect -611 357 -593 391
rect -559 357 -541 391
rect -483 357 -465 391
rect -431 357 -413 391
rect -355 357 -337 391
rect -303 357 -285 391
rect -227 357 -209 391
rect -175 357 -157 391
rect -99 357 -81 391
rect -47 357 -29 391
rect 29 357 47 391
rect 81 357 99 391
rect 157 357 175 391
rect 209 357 227 391
rect 285 357 303 391
rect 337 357 355 391
rect 413 357 431 391
rect 465 357 483 391
rect 541 357 559 391
rect 593 357 611 391
rect 669 357 687 391
rect 721 357 739 391
rect 797 357 815 391
rect 849 357 867 391
rect 925 357 943 391
rect 977 357 995 391
rect 1053 357 1071 391
rect 1105 357 1123 391
rect 1181 357 1199 391
rect 1233 357 1251 391
rect 1309 357 1327 391
rect 1361 357 1379 391
rect 1437 357 1455 391
rect 1489 357 1507 391
rect 1565 357 1583 391
rect 1617 357 1635 391
rect 1693 357 1711 391
rect 1745 357 1763 391
rect 1821 357 1839 391
rect 1873 357 1891 391
rect 1949 357 1967 391
rect 2001 357 2019 391
rect -2179 323 -2145 357
rect 2145 323 2179 357
rect -2179 255 -2145 289
rect -2179 187 -2145 221
rect -2179 119 -2145 153
rect -2179 51 -2145 85
rect -2179 -17 -2145 17
rect -2179 -85 -2145 -51
rect -2179 -153 -2145 -119
rect -2179 -221 -2145 -187
rect -2179 -289 -2145 -255
rect -2179 -357 -2145 -323
rect -2065 292 -2031 323
rect -2065 224 -2031 240
rect -2065 156 -2031 168
rect -2065 88 -2031 96
rect -2065 20 -2031 24
rect -2065 -86 -2031 -82
rect -2065 -158 -2031 -150
rect -2065 -230 -2031 -218
rect -2065 -302 -2031 -286
rect -2065 -385 -2031 -354
rect -1937 292 -1903 323
rect -1937 224 -1903 240
rect -1937 156 -1903 168
rect -1937 88 -1903 96
rect -1937 20 -1903 24
rect -1937 -86 -1903 -82
rect -1937 -158 -1903 -150
rect -1937 -230 -1903 -218
rect -1937 -302 -1903 -286
rect -1937 -385 -1903 -354
rect -1809 292 -1775 323
rect -1809 224 -1775 240
rect -1809 156 -1775 168
rect -1809 88 -1775 96
rect -1809 20 -1775 24
rect -1809 -86 -1775 -82
rect -1809 -158 -1775 -150
rect -1809 -230 -1775 -218
rect -1809 -302 -1775 -286
rect -1809 -385 -1775 -354
rect -1681 292 -1647 323
rect -1681 224 -1647 240
rect -1681 156 -1647 168
rect -1681 88 -1647 96
rect -1681 20 -1647 24
rect -1681 -86 -1647 -82
rect -1681 -158 -1647 -150
rect -1681 -230 -1647 -218
rect -1681 -302 -1647 -286
rect -1681 -385 -1647 -354
rect -1553 292 -1519 323
rect -1553 224 -1519 240
rect -1553 156 -1519 168
rect -1553 88 -1519 96
rect -1553 20 -1519 24
rect -1553 -86 -1519 -82
rect -1553 -158 -1519 -150
rect -1553 -230 -1519 -218
rect -1553 -302 -1519 -286
rect -1553 -385 -1519 -354
rect -1425 292 -1391 323
rect -1425 224 -1391 240
rect -1425 156 -1391 168
rect -1425 88 -1391 96
rect -1425 20 -1391 24
rect -1425 -86 -1391 -82
rect -1425 -158 -1391 -150
rect -1425 -230 -1391 -218
rect -1425 -302 -1391 -286
rect -1425 -385 -1391 -354
rect -1297 292 -1263 323
rect -1297 224 -1263 240
rect -1297 156 -1263 168
rect -1297 88 -1263 96
rect -1297 20 -1263 24
rect -1297 -86 -1263 -82
rect -1297 -158 -1263 -150
rect -1297 -230 -1263 -218
rect -1297 -302 -1263 -286
rect -1297 -385 -1263 -354
rect -1169 292 -1135 323
rect -1169 224 -1135 240
rect -1169 156 -1135 168
rect -1169 88 -1135 96
rect -1169 20 -1135 24
rect -1169 -86 -1135 -82
rect -1169 -158 -1135 -150
rect -1169 -230 -1135 -218
rect -1169 -302 -1135 -286
rect -1169 -385 -1135 -354
rect -1041 292 -1007 323
rect -1041 224 -1007 240
rect -1041 156 -1007 168
rect -1041 88 -1007 96
rect -1041 20 -1007 24
rect -1041 -86 -1007 -82
rect -1041 -158 -1007 -150
rect -1041 -230 -1007 -218
rect -1041 -302 -1007 -286
rect -1041 -385 -1007 -354
rect -913 292 -879 323
rect -913 224 -879 240
rect -913 156 -879 168
rect -913 88 -879 96
rect -913 20 -879 24
rect -913 -86 -879 -82
rect -913 -158 -879 -150
rect -913 -230 -879 -218
rect -913 -302 -879 -286
rect -913 -385 -879 -354
rect -785 292 -751 323
rect -785 224 -751 240
rect -785 156 -751 168
rect -785 88 -751 96
rect -785 20 -751 24
rect -785 -86 -751 -82
rect -785 -158 -751 -150
rect -785 -230 -751 -218
rect -785 -302 -751 -286
rect -785 -385 -751 -354
rect -657 292 -623 323
rect -657 224 -623 240
rect -657 156 -623 168
rect -657 88 -623 96
rect -657 20 -623 24
rect -657 -86 -623 -82
rect -657 -158 -623 -150
rect -657 -230 -623 -218
rect -657 -302 -623 -286
rect -657 -385 -623 -354
rect -529 292 -495 323
rect -529 224 -495 240
rect -529 156 -495 168
rect -529 88 -495 96
rect -529 20 -495 24
rect -529 -86 -495 -82
rect -529 -158 -495 -150
rect -529 -230 -495 -218
rect -529 -302 -495 -286
rect -529 -385 -495 -354
rect -401 292 -367 323
rect -401 224 -367 240
rect -401 156 -367 168
rect -401 88 -367 96
rect -401 20 -367 24
rect -401 -86 -367 -82
rect -401 -158 -367 -150
rect -401 -230 -367 -218
rect -401 -302 -367 -286
rect -401 -385 -367 -354
rect -273 292 -239 323
rect -273 224 -239 240
rect -273 156 -239 168
rect -273 88 -239 96
rect -273 20 -239 24
rect -273 -86 -239 -82
rect -273 -158 -239 -150
rect -273 -230 -239 -218
rect -273 -302 -239 -286
rect -273 -385 -239 -354
rect -145 292 -111 323
rect -145 224 -111 240
rect -145 156 -111 168
rect -145 88 -111 96
rect -145 20 -111 24
rect -145 -86 -111 -82
rect -145 -158 -111 -150
rect -145 -230 -111 -218
rect -145 -302 -111 -286
rect -145 -385 -111 -354
rect -17 292 17 323
rect -17 224 17 240
rect -17 156 17 168
rect -17 88 17 96
rect -17 20 17 24
rect -17 -86 17 -82
rect -17 -158 17 -150
rect -17 -230 17 -218
rect -17 -302 17 -286
rect -17 -385 17 -354
rect 111 292 145 323
rect 111 224 145 240
rect 111 156 145 168
rect 111 88 145 96
rect 111 20 145 24
rect 111 -86 145 -82
rect 111 -158 145 -150
rect 111 -230 145 -218
rect 111 -302 145 -286
rect 111 -385 145 -354
rect 239 292 273 323
rect 239 224 273 240
rect 239 156 273 168
rect 239 88 273 96
rect 239 20 273 24
rect 239 -86 273 -82
rect 239 -158 273 -150
rect 239 -230 273 -218
rect 239 -302 273 -286
rect 239 -385 273 -354
rect 367 292 401 323
rect 367 224 401 240
rect 367 156 401 168
rect 367 88 401 96
rect 367 20 401 24
rect 367 -86 401 -82
rect 367 -158 401 -150
rect 367 -230 401 -218
rect 367 -302 401 -286
rect 367 -385 401 -354
rect 495 292 529 323
rect 495 224 529 240
rect 495 156 529 168
rect 495 88 529 96
rect 495 20 529 24
rect 495 -86 529 -82
rect 495 -158 529 -150
rect 495 -230 529 -218
rect 495 -302 529 -286
rect 495 -385 529 -354
rect 623 292 657 323
rect 623 224 657 240
rect 623 156 657 168
rect 623 88 657 96
rect 623 20 657 24
rect 623 -86 657 -82
rect 623 -158 657 -150
rect 623 -230 657 -218
rect 623 -302 657 -286
rect 623 -385 657 -354
rect 751 292 785 323
rect 751 224 785 240
rect 751 156 785 168
rect 751 88 785 96
rect 751 20 785 24
rect 751 -86 785 -82
rect 751 -158 785 -150
rect 751 -230 785 -218
rect 751 -302 785 -286
rect 751 -385 785 -354
rect 879 292 913 323
rect 879 224 913 240
rect 879 156 913 168
rect 879 88 913 96
rect 879 20 913 24
rect 879 -86 913 -82
rect 879 -158 913 -150
rect 879 -230 913 -218
rect 879 -302 913 -286
rect 879 -385 913 -354
rect 1007 292 1041 323
rect 1007 224 1041 240
rect 1007 156 1041 168
rect 1007 88 1041 96
rect 1007 20 1041 24
rect 1007 -86 1041 -82
rect 1007 -158 1041 -150
rect 1007 -230 1041 -218
rect 1007 -302 1041 -286
rect 1007 -385 1041 -354
rect 1135 292 1169 323
rect 1135 224 1169 240
rect 1135 156 1169 168
rect 1135 88 1169 96
rect 1135 20 1169 24
rect 1135 -86 1169 -82
rect 1135 -158 1169 -150
rect 1135 -230 1169 -218
rect 1135 -302 1169 -286
rect 1135 -385 1169 -354
rect 1263 292 1297 323
rect 1263 224 1297 240
rect 1263 156 1297 168
rect 1263 88 1297 96
rect 1263 20 1297 24
rect 1263 -86 1297 -82
rect 1263 -158 1297 -150
rect 1263 -230 1297 -218
rect 1263 -302 1297 -286
rect 1263 -385 1297 -354
rect 1391 292 1425 323
rect 1391 224 1425 240
rect 1391 156 1425 168
rect 1391 88 1425 96
rect 1391 20 1425 24
rect 1391 -86 1425 -82
rect 1391 -158 1425 -150
rect 1391 -230 1425 -218
rect 1391 -302 1425 -286
rect 1391 -385 1425 -354
rect 1519 292 1553 323
rect 1519 224 1553 240
rect 1519 156 1553 168
rect 1519 88 1553 96
rect 1519 20 1553 24
rect 1519 -86 1553 -82
rect 1519 -158 1553 -150
rect 1519 -230 1553 -218
rect 1519 -302 1553 -286
rect 1519 -385 1553 -354
rect 1647 292 1681 323
rect 1647 224 1681 240
rect 1647 156 1681 168
rect 1647 88 1681 96
rect 1647 20 1681 24
rect 1647 -86 1681 -82
rect 1647 -158 1681 -150
rect 1647 -230 1681 -218
rect 1647 -302 1681 -286
rect 1647 -385 1681 -354
rect 1775 292 1809 323
rect 1775 224 1809 240
rect 1775 156 1809 168
rect 1775 88 1809 96
rect 1775 20 1809 24
rect 1775 -86 1809 -82
rect 1775 -158 1809 -150
rect 1775 -230 1809 -218
rect 1775 -302 1809 -286
rect 1775 -385 1809 -354
rect 1903 292 1937 323
rect 1903 224 1937 240
rect 1903 156 1937 168
rect 1903 88 1937 96
rect 1903 20 1937 24
rect 1903 -86 1937 -82
rect 1903 -158 1937 -150
rect 1903 -230 1937 -218
rect 1903 -302 1937 -286
rect 1903 -385 1937 -354
rect 2031 292 2065 323
rect 2031 224 2065 240
rect 2031 156 2065 168
rect 2031 88 2065 96
rect 2031 20 2065 24
rect 2031 -86 2065 -82
rect 2031 -158 2065 -150
rect 2031 -230 2065 -218
rect 2031 -302 2065 -286
rect 2031 -385 2065 -354
rect 2145 255 2179 289
rect 2145 187 2179 221
rect 2145 119 2179 153
rect 2145 51 2179 85
rect 2145 -17 2179 17
rect 2145 -85 2179 -51
rect 2145 -153 2179 -119
rect 2145 -221 2179 -187
rect 2145 -289 2179 -255
rect 2145 -357 2179 -323
rect -2179 -459 -2145 -391
rect 2145 -459 2179 -391
rect -2179 -493 -2057 -459
rect -2023 -493 -1989 -459
rect -1955 -493 -1921 -459
rect -1887 -493 -1853 -459
rect -1819 -493 -1785 -459
rect -1751 -493 -1717 -459
rect -1683 -493 -1649 -459
rect -1615 -493 -1581 -459
rect -1547 -493 -1513 -459
rect -1479 -493 -1445 -459
rect -1411 -493 -1377 -459
rect -1343 -493 -1309 -459
rect -1275 -493 -1241 -459
rect -1207 -493 -1173 -459
rect -1139 -493 -1105 -459
rect -1071 -493 -1037 -459
rect -1003 -493 -969 -459
rect -935 -493 -901 -459
rect -867 -493 -833 -459
rect -799 -493 -765 -459
rect -731 -493 -697 -459
rect -663 -493 -629 -459
rect -595 -493 -561 -459
rect -527 -493 -493 -459
rect -459 -493 -425 -459
rect -391 -493 -357 -459
rect -323 -493 -289 -459
rect -255 -493 -221 -459
rect -187 -493 -153 -459
rect -119 -493 -85 -459
rect -51 -493 -17 -459
rect 17 -493 51 -459
rect 85 -493 119 -459
rect 153 -493 187 -459
rect 221 -493 255 -459
rect 289 -493 323 -459
rect 357 -493 391 -459
rect 425 -493 459 -459
rect 493 -493 527 -459
rect 561 -493 595 -459
rect 629 -493 663 -459
rect 697 -493 731 -459
rect 765 -493 799 -459
rect 833 -493 867 -459
rect 901 -493 935 -459
rect 969 -493 1003 -459
rect 1037 -493 1071 -459
rect 1105 -493 1139 -459
rect 1173 -493 1207 -459
rect 1241 -493 1275 -459
rect 1309 -493 1343 -459
rect 1377 -493 1411 -459
rect 1445 -493 1479 -459
rect 1513 -493 1547 -459
rect 1581 -493 1615 -459
rect 1649 -493 1683 -459
rect 1717 -493 1751 -459
rect 1785 -493 1819 -459
rect 1853 -493 1887 -459
rect 1921 -493 1955 -459
rect 1989 -493 2023 -459
rect 2057 -493 2179 -459
<< viali >>
rect -2001 357 -1967 391
rect -1873 357 -1839 391
rect -1745 357 -1711 391
rect -1617 357 -1583 391
rect -1489 357 -1455 391
rect -1361 357 -1327 391
rect -1233 357 -1199 391
rect -1105 357 -1071 391
rect -977 357 -943 391
rect -849 357 -815 391
rect -721 357 -687 391
rect -593 357 -559 391
rect -465 357 -431 391
rect -337 357 -303 391
rect -209 357 -175 391
rect -81 357 -47 391
rect 47 357 81 391
rect 175 357 209 391
rect 303 357 337 391
rect 431 357 465 391
rect 559 357 593 391
rect 687 357 721 391
rect 815 357 849 391
rect 943 357 977 391
rect 1071 357 1105 391
rect 1199 357 1233 391
rect 1327 357 1361 391
rect 1455 357 1489 391
rect 1583 357 1617 391
rect 1711 357 1745 391
rect 1839 357 1873 391
rect 1967 357 2001 391
rect -2065 258 -2031 274
rect -2065 240 -2031 258
rect -2065 190 -2031 202
rect -2065 168 -2031 190
rect -2065 122 -2031 130
rect -2065 96 -2031 122
rect -2065 54 -2031 58
rect -2065 24 -2031 54
rect -2065 -48 -2031 -14
rect -2065 -116 -2031 -86
rect -2065 -120 -2031 -116
rect -2065 -184 -2031 -158
rect -2065 -192 -2031 -184
rect -2065 -252 -2031 -230
rect -2065 -264 -2031 -252
rect -2065 -320 -2031 -302
rect -2065 -336 -2031 -320
rect -1937 258 -1903 274
rect -1937 240 -1903 258
rect -1937 190 -1903 202
rect -1937 168 -1903 190
rect -1937 122 -1903 130
rect -1937 96 -1903 122
rect -1937 54 -1903 58
rect -1937 24 -1903 54
rect -1937 -48 -1903 -14
rect -1937 -116 -1903 -86
rect -1937 -120 -1903 -116
rect -1937 -184 -1903 -158
rect -1937 -192 -1903 -184
rect -1937 -252 -1903 -230
rect -1937 -264 -1903 -252
rect -1937 -320 -1903 -302
rect -1937 -336 -1903 -320
rect -1809 258 -1775 274
rect -1809 240 -1775 258
rect -1809 190 -1775 202
rect -1809 168 -1775 190
rect -1809 122 -1775 130
rect -1809 96 -1775 122
rect -1809 54 -1775 58
rect -1809 24 -1775 54
rect -1809 -48 -1775 -14
rect -1809 -116 -1775 -86
rect -1809 -120 -1775 -116
rect -1809 -184 -1775 -158
rect -1809 -192 -1775 -184
rect -1809 -252 -1775 -230
rect -1809 -264 -1775 -252
rect -1809 -320 -1775 -302
rect -1809 -336 -1775 -320
rect -1681 258 -1647 274
rect -1681 240 -1647 258
rect -1681 190 -1647 202
rect -1681 168 -1647 190
rect -1681 122 -1647 130
rect -1681 96 -1647 122
rect -1681 54 -1647 58
rect -1681 24 -1647 54
rect -1681 -48 -1647 -14
rect -1681 -116 -1647 -86
rect -1681 -120 -1647 -116
rect -1681 -184 -1647 -158
rect -1681 -192 -1647 -184
rect -1681 -252 -1647 -230
rect -1681 -264 -1647 -252
rect -1681 -320 -1647 -302
rect -1681 -336 -1647 -320
rect -1553 258 -1519 274
rect -1553 240 -1519 258
rect -1553 190 -1519 202
rect -1553 168 -1519 190
rect -1553 122 -1519 130
rect -1553 96 -1519 122
rect -1553 54 -1519 58
rect -1553 24 -1519 54
rect -1553 -48 -1519 -14
rect -1553 -116 -1519 -86
rect -1553 -120 -1519 -116
rect -1553 -184 -1519 -158
rect -1553 -192 -1519 -184
rect -1553 -252 -1519 -230
rect -1553 -264 -1519 -252
rect -1553 -320 -1519 -302
rect -1553 -336 -1519 -320
rect -1425 258 -1391 274
rect -1425 240 -1391 258
rect -1425 190 -1391 202
rect -1425 168 -1391 190
rect -1425 122 -1391 130
rect -1425 96 -1391 122
rect -1425 54 -1391 58
rect -1425 24 -1391 54
rect -1425 -48 -1391 -14
rect -1425 -116 -1391 -86
rect -1425 -120 -1391 -116
rect -1425 -184 -1391 -158
rect -1425 -192 -1391 -184
rect -1425 -252 -1391 -230
rect -1425 -264 -1391 -252
rect -1425 -320 -1391 -302
rect -1425 -336 -1391 -320
rect -1297 258 -1263 274
rect -1297 240 -1263 258
rect -1297 190 -1263 202
rect -1297 168 -1263 190
rect -1297 122 -1263 130
rect -1297 96 -1263 122
rect -1297 54 -1263 58
rect -1297 24 -1263 54
rect -1297 -48 -1263 -14
rect -1297 -116 -1263 -86
rect -1297 -120 -1263 -116
rect -1297 -184 -1263 -158
rect -1297 -192 -1263 -184
rect -1297 -252 -1263 -230
rect -1297 -264 -1263 -252
rect -1297 -320 -1263 -302
rect -1297 -336 -1263 -320
rect -1169 258 -1135 274
rect -1169 240 -1135 258
rect -1169 190 -1135 202
rect -1169 168 -1135 190
rect -1169 122 -1135 130
rect -1169 96 -1135 122
rect -1169 54 -1135 58
rect -1169 24 -1135 54
rect -1169 -48 -1135 -14
rect -1169 -116 -1135 -86
rect -1169 -120 -1135 -116
rect -1169 -184 -1135 -158
rect -1169 -192 -1135 -184
rect -1169 -252 -1135 -230
rect -1169 -264 -1135 -252
rect -1169 -320 -1135 -302
rect -1169 -336 -1135 -320
rect -1041 258 -1007 274
rect -1041 240 -1007 258
rect -1041 190 -1007 202
rect -1041 168 -1007 190
rect -1041 122 -1007 130
rect -1041 96 -1007 122
rect -1041 54 -1007 58
rect -1041 24 -1007 54
rect -1041 -48 -1007 -14
rect -1041 -116 -1007 -86
rect -1041 -120 -1007 -116
rect -1041 -184 -1007 -158
rect -1041 -192 -1007 -184
rect -1041 -252 -1007 -230
rect -1041 -264 -1007 -252
rect -1041 -320 -1007 -302
rect -1041 -336 -1007 -320
rect -913 258 -879 274
rect -913 240 -879 258
rect -913 190 -879 202
rect -913 168 -879 190
rect -913 122 -879 130
rect -913 96 -879 122
rect -913 54 -879 58
rect -913 24 -879 54
rect -913 -48 -879 -14
rect -913 -116 -879 -86
rect -913 -120 -879 -116
rect -913 -184 -879 -158
rect -913 -192 -879 -184
rect -913 -252 -879 -230
rect -913 -264 -879 -252
rect -913 -320 -879 -302
rect -913 -336 -879 -320
rect -785 258 -751 274
rect -785 240 -751 258
rect -785 190 -751 202
rect -785 168 -751 190
rect -785 122 -751 130
rect -785 96 -751 122
rect -785 54 -751 58
rect -785 24 -751 54
rect -785 -48 -751 -14
rect -785 -116 -751 -86
rect -785 -120 -751 -116
rect -785 -184 -751 -158
rect -785 -192 -751 -184
rect -785 -252 -751 -230
rect -785 -264 -751 -252
rect -785 -320 -751 -302
rect -785 -336 -751 -320
rect -657 258 -623 274
rect -657 240 -623 258
rect -657 190 -623 202
rect -657 168 -623 190
rect -657 122 -623 130
rect -657 96 -623 122
rect -657 54 -623 58
rect -657 24 -623 54
rect -657 -48 -623 -14
rect -657 -116 -623 -86
rect -657 -120 -623 -116
rect -657 -184 -623 -158
rect -657 -192 -623 -184
rect -657 -252 -623 -230
rect -657 -264 -623 -252
rect -657 -320 -623 -302
rect -657 -336 -623 -320
rect -529 258 -495 274
rect -529 240 -495 258
rect -529 190 -495 202
rect -529 168 -495 190
rect -529 122 -495 130
rect -529 96 -495 122
rect -529 54 -495 58
rect -529 24 -495 54
rect -529 -48 -495 -14
rect -529 -116 -495 -86
rect -529 -120 -495 -116
rect -529 -184 -495 -158
rect -529 -192 -495 -184
rect -529 -252 -495 -230
rect -529 -264 -495 -252
rect -529 -320 -495 -302
rect -529 -336 -495 -320
rect -401 258 -367 274
rect -401 240 -367 258
rect -401 190 -367 202
rect -401 168 -367 190
rect -401 122 -367 130
rect -401 96 -367 122
rect -401 54 -367 58
rect -401 24 -367 54
rect -401 -48 -367 -14
rect -401 -116 -367 -86
rect -401 -120 -367 -116
rect -401 -184 -367 -158
rect -401 -192 -367 -184
rect -401 -252 -367 -230
rect -401 -264 -367 -252
rect -401 -320 -367 -302
rect -401 -336 -367 -320
rect -273 258 -239 274
rect -273 240 -239 258
rect -273 190 -239 202
rect -273 168 -239 190
rect -273 122 -239 130
rect -273 96 -239 122
rect -273 54 -239 58
rect -273 24 -239 54
rect -273 -48 -239 -14
rect -273 -116 -239 -86
rect -273 -120 -239 -116
rect -273 -184 -239 -158
rect -273 -192 -239 -184
rect -273 -252 -239 -230
rect -273 -264 -239 -252
rect -273 -320 -239 -302
rect -273 -336 -239 -320
rect -145 258 -111 274
rect -145 240 -111 258
rect -145 190 -111 202
rect -145 168 -111 190
rect -145 122 -111 130
rect -145 96 -111 122
rect -145 54 -111 58
rect -145 24 -111 54
rect -145 -48 -111 -14
rect -145 -116 -111 -86
rect -145 -120 -111 -116
rect -145 -184 -111 -158
rect -145 -192 -111 -184
rect -145 -252 -111 -230
rect -145 -264 -111 -252
rect -145 -320 -111 -302
rect -145 -336 -111 -320
rect -17 258 17 274
rect -17 240 17 258
rect -17 190 17 202
rect -17 168 17 190
rect -17 122 17 130
rect -17 96 17 122
rect -17 54 17 58
rect -17 24 17 54
rect -17 -48 17 -14
rect -17 -116 17 -86
rect -17 -120 17 -116
rect -17 -184 17 -158
rect -17 -192 17 -184
rect -17 -252 17 -230
rect -17 -264 17 -252
rect -17 -320 17 -302
rect -17 -336 17 -320
rect 111 258 145 274
rect 111 240 145 258
rect 111 190 145 202
rect 111 168 145 190
rect 111 122 145 130
rect 111 96 145 122
rect 111 54 145 58
rect 111 24 145 54
rect 111 -48 145 -14
rect 111 -116 145 -86
rect 111 -120 145 -116
rect 111 -184 145 -158
rect 111 -192 145 -184
rect 111 -252 145 -230
rect 111 -264 145 -252
rect 111 -320 145 -302
rect 111 -336 145 -320
rect 239 258 273 274
rect 239 240 273 258
rect 239 190 273 202
rect 239 168 273 190
rect 239 122 273 130
rect 239 96 273 122
rect 239 54 273 58
rect 239 24 273 54
rect 239 -48 273 -14
rect 239 -116 273 -86
rect 239 -120 273 -116
rect 239 -184 273 -158
rect 239 -192 273 -184
rect 239 -252 273 -230
rect 239 -264 273 -252
rect 239 -320 273 -302
rect 239 -336 273 -320
rect 367 258 401 274
rect 367 240 401 258
rect 367 190 401 202
rect 367 168 401 190
rect 367 122 401 130
rect 367 96 401 122
rect 367 54 401 58
rect 367 24 401 54
rect 367 -48 401 -14
rect 367 -116 401 -86
rect 367 -120 401 -116
rect 367 -184 401 -158
rect 367 -192 401 -184
rect 367 -252 401 -230
rect 367 -264 401 -252
rect 367 -320 401 -302
rect 367 -336 401 -320
rect 495 258 529 274
rect 495 240 529 258
rect 495 190 529 202
rect 495 168 529 190
rect 495 122 529 130
rect 495 96 529 122
rect 495 54 529 58
rect 495 24 529 54
rect 495 -48 529 -14
rect 495 -116 529 -86
rect 495 -120 529 -116
rect 495 -184 529 -158
rect 495 -192 529 -184
rect 495 -252 529 -230
rect 495 -264 529 -252
rect 495 -320 529 -302
rect 495 -336 529 -320
rect 623 258 657 274
rect 623 240 657 258
rect 623 190 657 202
rect 623 168 657 190
rect 623 122 657 130
rect 623 96 657 122
rect 623 54 657 58
rect 623 24 657 54
rect 623 -48 657 -14
rect 623 -116 657 -86
rect 623 -120 657 -116
rect 623 -184 657 -158
rect 623 -192 657 -184
rect 623 -252 657 -230
rect 623 -264 657 -252
rect 623 -320 657 -302
rect 623 -336 657 -320
rect 751 258 785 274
rect 751 240 785 258
rect 751 190 785 202
rect 751 168 785 190
rect 751 122 785 130
rect 751 96 785 122
rect 751 54 785 58
rect 751 24 785 54
rect 751 -48 785 -14
rect 751 -116 785 -86
rect 751 -120 785 -116
rect 751 -184 785 -158
rect 751 -192 785 -184
rect 751 -252 785 -230
rect 751 -264 785 -252
rect 751 -320 785 -302
rect 751 -336 785 -320
rect 879 258 913 274
rect 879 240 913 258
rect 879 190 913 202
rect 879 168 913 190
rect 879 122 913 130
rect 879 96 913 122
rect 879 54 913 58
rect 879 24 913 54
rect 879 -48 913 -14
rect 879 -116 913 -86
rect 879 -120 913 -116
rect 879 -184 913 -158
rect 879 -192 913 -184
rect 879 -252 913 -230
rect 879 -264 913 -252
rect 879 -320 913 -302
rect 879 -336 913 -320
rect 1007 258 1041 274
rect 1007 240 1041 258
rect 1007 190 1041 202
rect 1007 168 1041 190
rect 1007 122 1041 130
rect 1007 96 1041 122
rect 1007 54 1041 58
rect 1007 24 1041 54
rect 1007 -48 1041 -14
rect 1007 -116 1041 -86
rect 1007 -120 1041 -116
rect 1007 -184 1041 -158
rect 1007 -192 1041 -184
rect 1007 -252 1041 -230
rect 1007 -264 1041 -252
rect 1007 -320 1041 -302
rect 1007 -336 1041 -320
rect 1135 258 1169 274
rect 1135 240 1169 258
rect 1135 190 1169 202
rect 1135 168 1169 190
rect 1135 122 1169 130
rect 1135 96 1169 122
rect 1135 54 1169 58
rect 1135 24 1169 54
rect 1135 -48 1169 -14
rect 1135 -116 1169 -86
rect 1135 -120 1169 -116
rect 1135 -184 1169 -158
rect 1135 -192 1169 -184
rect 1135 -252 1169 -230
rect 1135 -264 1169 -252
rect 1135 -320 1169 -302
rect 1135 -336 1169 -320
rect 1263 258 1297 274
rect 1263 240 1297 258
rect 1263 190 1297 202
rect 1263 168 1297 190
rect 1263 122 1297 130
rect 1263 96 1297 122
rect 1263 54 1297 58
rect 1263 24 1297 54
rect 1263 -48 1297 -14
rect 1263 -116 1297 -86
rect 1263 -120 1297 -116
rect 1263 -184 1297 -158
rect 1263 -192 1297 -184
rect 1263 -252 1297 -230
rect 1263 -264 1297 -252
rect 1263 -320 1297 -302
rect 1263 -336 1297 -320
rect 1391 258 1425 274
rect 1391 240 1425 258
rect 1391 190 1425 202
rect 1391 168 1425 190
rect 1391 122 1425 130
rect 1391 96 1425 122
rect 1391 54 1425 58
rect 1391 24 1425 54
rect 1391 -48 1425 -14
rect 1391 -116 1425 -86
rect 1391 -120 1425 -116
rect 1391 -184 1425 -158
rect 1391 -192 1425 -184
rect 1391 -252 1425 -230
rect 1391 -264 1425 -252
rect 1391 -320 1425 -302
rect 1391 -336 1425 -320
rect 1519 258 1553 274
rect 1519 240 1553 258
rect 1519 190 1553 202
rect 1519 168 1553 190
rect 1519 122 1553 130
rect 1519 96 1553 122
rect 1519 54 1553 58
rect 1519 24 1553 54
rect 1519 -48 1553 -14
rect 1519 -116 1553 -86
rect 1519 -120 1553 -116
rect 1519 -184 1553 -158
rect 1519 -192 1553 -184
rect 1519 -252 1553 -230
rect 1519 -264 1553 -252
rect 1519 -320 1553 -302
rect 1519 -336 1553 -320
rect 1647 258 1681 274
rect 1647 240 1681 258
rect 1647 190 1681 202
rect 1647 168 1681 190
rect 1647 122 1681 130
rect 1647 96 1681 122
rect 1647 54 1681 58
rect 1647 24 1681 54
rect 1647 -48 1681 -14
rect 1647 -116 1681 -86
rect 1647 -120 1681 -116
rect 1647 -184 1681 -158
rect 1647 -192 1681 -184
rect 1647 -252 1681 -230
rect 1647 -264 1681 -252
rect 1647 -320 1681 -302
rect 1647 -336 1681 -320
rect 1775 258 1809 274
rect 1775 240 1809 258
rect 1775 190 1809 202
rect 1775 168 1809 190
rect 1775 122 1809 130
rect 1775 96 1809 122
rect 1775 54 1809 58
rect 1775 24 1809 54
rect 1775 -48 1809 -14
rect 1775 -116 1809 -86
rect 1775 -120 1809 -116
rect 1775 -184 1809 -158
rect 1775 -192 1809 -184
rect 1775 -252 1809 -230
rect 1775 -264 1809 -252
rect 1775 -320 1809 -302
rect 1775 -336 1809 -320
rect 1903 258 1937 274
rect 1903 240 1937 258
rect 1903 190 1937 202
rect 1903 168 1937 190
rect 1903 122 1937 130
rect 1903 96 1937 122
rect 1903 54 1937 58
rect 1903 24 1937 54
rect 1903 -48 1937 -14
rect 1903 -116 1937 -86
rect 1903 -120 1937 -116
rect 1903 -184 1937 -158
rect 1903 -192 1937 -184
rect 1903 -252 1937 -230
rect 1903 -264 1937 -252
rect 1903 -320 1937 -302
rect 1903 -336 1937 -320
rect 2031 258 2065 274
rect 2031 240 2065 258
rect 2031 190 2065 202
rect 2031 168 2065 190
rect 2031 122 2065 130
rect 2031 96 2065 122
rect 2031 54 2065 58
rect 2031 24 2065 54
rect 2031 -48 2065 -14
rect 2031 -116 2065 -86
rect 2031 -120 2065 -116
rect 2031 -184 2065 -158
rect 2031 -192 2065 -184
rect 2031 -252 2065 -230
rect 2031 -264 2065 -252
rect 2031 -320 2065 -302
rect 2031 -336 2065 -320
<< metal1 >>
rect -2015 391 -1953 397
rect -2015 357 -2001 391
rect -1967 357 -1953 391
rect -2015 351 -1953 357
rect -1887 391 -1825 397
rect -1887 357 -1873 391
rect -1839 357 -1825 391
rect -1887 351 -1825 357
rect -1759 391 -1697 397
rect -1759 357 -1745 391
rect -1711 357 -1697 391
rect -1759 351 -1697 357
rect -1631 391 -1569 397
rect -1631 357 -1617 391
rect -1583 357 -1569 391
rect -1631 351 -1569 357
rect -1503 391 -1441 397
rect -1503 357 -1489 391
rect -1455 357 -1441 391
rect -1503 351 -1441 357
rect -1375 391 -1313 397
rect -1375 357 -1361 391
rect -1327 357 -1313 391
rect -1375 351 -1313 357
rect -1247 391 -1185 397
rect -1247 357 -1233 391
rect -1199 357 -1185 391
rect -1247 351 -1185 357
rect -1119 391 -1057 397
rect -1119 357 -1105 391
rect -1071 357 -1057 391
rect -1119 351 -1057 357
rect -991 391 -929 397
rect -991 357 -977 391
rect -943 357 -929 391
rect -991 351 -929 357
rect -863 391 -801 397
rect -863 357 -849 391
rect -815 357 -801 391
rect -863 351 -801 357
rect -735 391 -673 397
rect -735 357 -721 391
rect -687 357 -673 391
rect -735 351 -673 357
rect -607 391 -545 397
rect -607 357 -593 391
rect -559 357 -545 391
rect -607 351 -545 357
rect -479 391 -417 397
rect -479 357 -465 391
rect -431 357 -417 391
rect -479 351 -417 357
rect -351 391 -289 397
rect -351 357 -337 391
rect -303 357 -289 391
rect -351 351 -289 357
rect -223 391 -161 397
rect -223 357 -209 391
rect -175 357 -161 391
rect -223 351 -161 357
rect -95 391 -33 397
rect -95 357 -81 391
rect -47 357 -33 391
rect -95 351 -33 357
rect 33 391 95 397
rect 33 357 47 391
rect 81 357 95 391
rect 33 351 95 357
rect 161 391 223 397
rect 161 357 175 391
rect 209 357 223 391
rect 161 351 223 357
rect 289 391 351 397
rect 289 357 303 391
rect 337 357 351 391
rect 289 351 351 357
rect 417 391 479 397
rect 417 357 431 391
rect 465 357 479 391
rect 417 351 479 357
rect 545 391 607 397
rect 545 357 559 391
rect 593 357 607 391
rect 545 351 607 357
rect 673 391 735 397
rect 673 357 687 391
rect 721 357 735 391
rect 673 351 735 357
rect 801 391 863 397
rect 801 357 815 391
rect 849 357 863 391
rect 801 351 863 357
rect 929 391 991 397
rect 929 357 943 391
rect 977 357 991 391
rect 929 351 991 357
rect 1057 391 1119 397
rect 1057 357 1071 391
rect 1105 357 1119 391
rect 1057 351 1119 357
rect 1185 391 1247 397
rect 1185 357 1199 391
rect 1233 357 1247 391
rect 1185 351 1247 357
rect 1313 391 1375 397
rect 1313 357 1327 391
rect 1361 357 1375 391
rect 1313 351 1375 357
rect 1441 391 1503 397
rect 1441 357 1455 391
rect 1489 357 1503 391
rect 1441 351 1503 357
rect 1569 391 1631 397
rect 1569 357 1583 391
rect 1617 357 1631 391
rect 1569 351 1631 357
rect 1697 391 1759 397
rect 1697 357 1711 391
rect 1745 357 1759 391
rect 1697 351 1759 357
rect 1825 391 1887 397
rect 1825 357 1839 391
rect 1873 357 1887 391
rect 1825 351 1887 357
rect 1953 391 2015 397
rect 1953 357 1967 391
rect 2001 357 2015 391
rect 1953 351 2015 357
rect -2071 274 -2025 319
rect -2071 240 -2065 274
rect -2031 240 -2025 274
rect -2071 202 -2025 240
rect -2071 168 -2065 202
rect -2031 168 -2025 202
rect -2071 130 -2025 168
rect -2071 96 -2065 130
rect -2031 96 -2025 130
rect -2071 58 -2025 96
rect -2071 24 -2065 58
rect -2031 24 -2025 58
rect -2071 -14 -2025 24
rect -2071 -48 -2065 -14
rect -2031 -48 -2025 -14
rect -2071 -86 -2025 -48
rect -2071 -120 -2065 -86
rect -2031 -120 -2025 -86
rect -2071 -158 -2025 -120
rect -2071 -192 -2065 -158
rect -2031 -192 -2025 -158
rect -2071 -230 -2025 -192
rect -2071 -264 -2065 -230
rect -2031 -264 -2025 -230
rect -2071 -302 -2025 -264
rect -2071 -336 -2065 -302
rect -2031 -336 -2025 -302
rect -2071 -381 -2025 -336
rect -1943 274 -1897 319
rect -1943 240 -1937 274
rect -1903 240 -1897 274
rect -1943 202 -1897 240
rect -1943 168 -1937 202
rect -1903 168 -1897 202
rect -1943 130 -1897 168
rect -1943 96 -1937 130
rect -1903 96 -1897 130
rect -1943 58 -1897 96
rect -1943 24 -1937 58
rect -1903 24 -1897 58
rect -1943 -14 -1897 24
rect -1943 -48 -1937 -14
rect -1903 -48 -1897 -14
rect -1943 -86 -1897 -48
rect -1943 -120 -1937 -86
rect -1903 -120 -1897 -86
rect -1943 -158 -1897 -120
rect -1943 -192 -1937 -158
rect -1903 -192 -1897 -158
rect -1943 -230 -1897 -192
rect -1943 -264 -1937 -230
rect -1903 -264 -1897 -230
rect -1943 -302 -1897 -264
rect -1943 -336 -1937 -302
rect -1903 -336 -1897 -302
rect -1943 -381 -1897 -336
rect -1815 274 -1769 319
rect -1815 240 -1809 274
rect -1775 240 -1769 274
rect -1815 202 -1769 240
rect -1815 168 -1809 202
rect -1775 168 -1769 202
rect -1815 130 -1769 168
rect -1815 96 -1809 130
rect -1775 96 -1769 130
rect -1815 58 -1769 96
rect -1815 24 -1809 58
rect -1775 24 -1769 58
rect -1815 -14 -1769 24
rect -1815 -48 -1809 -14
rect -1775 -48 -1769 -14
rect -1815 -86 -1769 -48
rect -1815 -120 -1809 -86
rect -1775 -120 -1769 -86
rect -1815 -158 -1769 -120
rect -1815 -192 -1809 -158
rect -1775 -192 -1769 -158
rect -1815 -230 -1769 -192
rect -1815 -264 -1809 -230
rect -1775 -264 -1769 -230
rect -1815 -302 -1769 -264
rect -1815 -336 -1809 -302
rect -1775 -336 -1769 -302
rect -1815 -381 -1769 -336
rect -1687 274 -1641 319
rect -1687 240 -1681 274
rect -1647 240 -1641 274
rect -1687 202 -1641 240
rect -1687 168 -1681 202
rect -1647 168 -1641 202
rect -1687 130 -1641 168
rect -1687 96 -1681 130
rect -1647 96 -1641 130
rect -1687 58 -1641 96
rect -1687 24 -1681 58
rect -1647 24 -1641 58
rect -1687 -14 -1641 24
rect -1687 -48 -1681 -14
rect -1647 -48 -1641 -14
rect -1687 -86 -1641 -48
rect -1687 -120 -1681 -86
rect -1647 -120 -1641 -86
rect -1687 -158 -1641 -120
rect -1687 -192 -1681 -158
rect -1647 -192 -1641 -158
rect -1687 -230 -1641 -192
rect -1687 -264 -1681 -230
rect -1647 -264 -1641 -230
rect -1687 -302 -1641 -264
rect -1687 -336 -1681 -302
rect -1647 -336 -1641 -302
rect -1687 -381 -1641 -336
rect -1559 274 -1513 319
rect -1559 240 -1553 274
rect -1519 240 -1513 274
rect -1559 202 -1513 240
rect -1559 168 -1553 202
rect -1519 168 -1513 202
rect -1559 130 -1513 168
rect -1559 96 -1553 130
rect -1519 96 -1513 130
rect -1559 58 -1513 96
rect -1559 24 -1553 58
rect -1519 24 -1513 58
rect -1559 -14 -1513 24
rect -1559 -48 -1553 -14
rect -1519 -48 -1513 -14
rect -1559 -86 -1513 -48
rect -1559 -120 -1553 -86
rect -1519 -120 -1513 -86
rect -1559 -158 -1513 -120
rect -1559 -192 -1553 -158
rect -1519 -192 -1513 -158
rect -1559 -230 -1513 -192
rect -1559 -264 -1553 -230
rect -1519 -264 -1513 -230
rect -1559 -302 -1513 -264
rect -1559 -336 -1553 -302
rect -1519 -336 -1513 -302
rect -1559 -381 -1513 -336
rect -1431 274 -1385 319
rect -1431 240 -1425 274
rect -1391 240 -1385 274
rect -1431 202 -1385 240
rect -1431 168 -1425 202
rect -1391 168 -1385 202
rect -1431 130 -1385 168
rect -1431 96 -1425 130
rect -1391 96 -1385 130
rect -1431 58 -1385 96
rect -1431 24 -1425 58
rect -1391 24 -1385 58
rect -1431 -14 -1385 24
rect -1431 -48 -1425 -14
rect -1391 -48 -1385 -14
rect -1431 -86 -1385 -48
rect -1431 -120 -1425 -86
rect -1391 -120 -1385 -86
rect -1431 -158 -1385 -120
rect -1431 -192 -1425 -158
rect -1391 -192 -1385 -158
rect -1431 -230 -1385 -192
rect -1431 -264 -1425 -230
rect -1391 -264 -1385 -230
rect -1431 -302 -1385 -264
rect -1431 -336 -1425 -302
rect -1391 -336 -1385 -302
rect -1431 -381 -1385 -336
rect -1303 274 -1257 319
rect -1303 240 -1297 274
rect -1263 240 -1257 274
rect -1303 202 -1257 240
rect -1303 168 -1297 202
rect -1263 168 -1257 202
rect -1303 130 -1257 168
rect -1303 96 -1297 130
rect -1263 96 -1257 130
rect -1303 58 -1257 96
rect -1303 24 -1297 58
rect -1263 24 -1257 58
rect -1303 -14 -1257 24
rect -1303 -48 -1297 -14
rect -1263 -48 -1257 -14
rect -1303 -86 -1257 -48
rect -1303 -120 -1297 -86
rect -1263 -120 -1257 -86
rect -1303 -158 -1257 -120
rect -1303 -192 -1297 -158
rect -1263 -192 -1257 -158
rect -1303 -230 -1257 -192
rect -1303 -264 -1297 -230
rect -1263 -264 -1257 -230
rect -1303 -302 -1257 -264
rect -1303 -336 -1297 -302
rect -1263 -336 -1257 -302
rect -1303 -381 -1257 -336
rect -1175 274 -1129 319
rect -1175 240 -1169 274
rect -1135 240 -1129 274
rect -1175 202 -1129 240
rect -1175 168 -1169 202
rect -1135 168 -1129 202
rect -1175 130 -1129 168
rect -1175 96 -1169 130
rect -1135 96 -1129 130
rect -1175 58 -1129 96
rect -1175 24 -1169 58
rect -1135 24 -1129 58
rect -1175 -14 -1129 24
rect -1175 -48 -1169 -14
rect -1135 -48 -1129 -14
rect -1175 -86 -1129 -48
rect -1175 -120 -1169 -86
rect -1135 -120 -1129 -86
rect -1175 -158 -1129 -120
rect -1175 -192 -1169 -158
rect -1135 -192 -1129 -158
rect -1175 -230 -1129 -192
rect -1175 -264 -1169 -230
rect -1135 -264 -1129 -230
rect -1175 -302 -1129 -264
rect -1175 -336 -1169 -302
rect -1135 -336 -1129 -302
rect -1175 -381 -1129 -336
rect -1047 274 -1001 319
rect -1047 240 -1041 274
rect -1007 240 -1001 274
rect -1047 202 -1001 240
rect -1047 168 -1041 202
rect -1007 168 -1001 202
rect -1047 130 -1001 168
rect -1047 96 -1041 130
rect -1007 96 -1001 130
rect -1047 58 -1001 96
rect -1047 24 -1041 58
rect -1007 24 -1001 58
rect -1047 -14 -1001 24
rect -1047 -48 -1041 -14
rect -1007 -48 -1001 -14
rect -1047 -86 -1001 -48
rect -1047 -120 -1041 -86
rect -1007 -120 -1001 -86
rect -1047 -158 -1001 -120
rect -1047 -192 -1041 -158
rect -1007 -192 -1001 -158
rect -1047 -230 -1001 -192
rect -1047 -264 -1041 -230
rect -1007 -264 -1001 -230
rect -1047 -302 -1001 -264
rect -1047 -336 -1041 -302
rect -1007 -336 -1001 -302
rect -1047 -381 -1001 -336
rect -919 274 -873 319
rect -919 240 -913 274
rect -879 240 -873 274
rect -919 202 -873 240
rect -919 168 -913 202
rect -879 168 -873 202
rect -919 130 -873 168
rect -919 96 -913 130
rect -879 96 -873 130
rect -919 58 -873 96
rect -919 24 -913 58
rect -879 24 -873 58
rect -919 -14 -873 24
rect -919 -48 -913 -14
rect -879 -48 -873 -14
rect -919 -86 -873 -48
rect -919 -120 -913 -86
rect -879 -120 -873 -86
rect -919 -158 -873 -120
rect -919 -192 -913 -158
rect -879 -192 -873 -158
rect -919 -230 -873 -192
rect -919 -264 -913 -230
rect -879 -264 -873 -230
rect -919 -302 -873 -264
rect -919 -336 -913 -302
rect -879 -336 -873 -302
rect -919 -381 -873 -336
rect -791 274 -745 319
rect -791 240 -785 274
rect -751 240 -745 274
rect -791 202 -745 240
rect -791 168 -785 202
rect -751 168 -745 202
rect -791 130 -745 168
rect -791 96 -785 130
rect -751 96 -745 130
rect -791 58 -745 96
rect -791 24 -785 58
rect -751 24 -745 58
rect -791 -14 -745 24
rect -791 -48 -785 -14
rect -751 -48 -745 -14
rect -791 -86 -745 -48
rect -791 -120 -785 -86
rect -751 -120 -745 -86
rect -791 -158 -745 -120
rect -791 -192 -785 -158
rect -751 -192 -745 -158
rect -791 -230 -745 -192
rect -791 -264 -785 -230
rect -751 -264 -745 -230
rect -791 -302 -745 -264
rect -791 -336 -785 -302
rect -751 -336 -745 -302
rect -791 -381 -745 -336
rect -663 274 -617 319
rect -663 240 -657 274
rect -623 240 -617 274
rect -663 202 -617 240
rect -663 168 -657 202
rect -623 168 -617 202
rect -663 130 -617 168
rect -663 96 -657 130
rect -623 96 -617 130
rect -663 58 -617 96
rect -663 24 -657 58
rect -623 24 -617 58
rect -663 -14 -617 24
rect -663 -48 -657 -14
rect -623 -48 -617 -14
rect -663 -86 -617 -48
rect -663 -120 -657 -86
rect -623 -120 -617 -86
rect -663 -158 -617 -120
rect -663 -192 -657 -158
rect -623 -192 -617 -158
rect -663 -230 -617 -192
rect -663 -264 -657 -230
rect -623 -264 -617 -230
rect -663 -302 -617 -264
rect -663 -336 -657 -302
rect -623 -336 -617 -302
rect -663 -381 -617 -336
rect -535 274 -489 319
rect -535 240 -529 274
rect -495 240 -489 274
rect -535 202 -489 240
rect -535 168 -529 202
rect -495 168 -489 202
rect -535 130 -489 168
rect -535 96 -529 130
rect -495 96 -489 130
rect -535 58 -489 96
rect -535 24 -529 58
rect -495 24 -489 58
rect -535 -14 -489 24
rect -535 -48 -529 -14
rect -495 -48 -489 -14
rect -535 -86 -489 -48
rect -535 -120 -529 -86
rect -495 -120 -489 -86
rect -535 -158 -489 -120
rect -535 -192 -529 -158
rect -495 -192 -489 -158
rect -535 -230 -489 -192
rect -535 -264 -529 -230
rect -495 -264 -489 -230
rect -535 -302 -489 -264
rect -535 -336 -529 -302
rect -495 -336 -489 -302
rect -535 -381 -489 -336
rect -407 274 -361 319
rect -407 240 -401 274
rect -367 240 -361 274
rect -407 202 -361 240
rect -407 168 -401 202
rect -367 168 -361 202
rect -407 130 -361 168
rect -407 96 -401 130
rect -367 96 -361 130
rect -407 58 -361 96
rect -407 24 -401 58
rect -367 24 -361 58
rect -407 -14 -361 24
rect -407 -48 -401 -14
rect -367 -48 -361 -14
rect -407 -86 -361 -48
rect -407 -120 -401 -86
rect -367 -120 -361 -86
rect -407 -158 -361 -120
rect -407 -192 -401 -158
rect -367 -192 -361 -158
rect -407 -230 -361 -192
rect -407 -264 -401 -230
rect -367 -264 -361 -230
rect -407 -302 -361 -264
rect -407 -336 -401 -302
rect -367 -336 -361 -302
rect -407 -381 -361 -336
rect -279 274 -233 319
rect -279 240 -273 274
rect -239 240 -233 274
rect -279 202 -233 240
rect -279 168 -273 202
rect -239 168 -233 202
rect -279 130 -233 168
rect -279 96 -273 130
rect -239 96 -233 130
rect -279 58 -233 96
rect -279 24 -273 58
rect -239 24 -233 58
rect -279 -14 -233 24
rect -279 -48 -273 -14
rect -239 -48 -233 -14
rect -279 -86 -233 -48
rect -279 -120 -273 -86
rect -239 -120 -233 -86
rect -279 -158 -233 -120
rect -279 -192 -273 -158
rect -239 -192 -233 -158
rect -279 -230 -233 -192
rect -279 -264 -273 -230
rect -239 -264 -233 -230
rect -279 -302 -233 -264
rect -279 -336 -273 -302
rect -239 -336 -233 -302
rect -279 -381 -233 -336
rect -151 274 -105 319
rect -151 240 -145 274
rect -111 240 -105 274
rect -151 202 -105 240
rect -151 168 -145 202
rect -111 168 -105 202
rect -151 130 -105 168
rect -151 96 -145 130
rect -111 96 -105 130
rect -151 58 -105 96
rect -151 24 -145 58
rect -111 24 -105 58
rect -151 -14 -105 24
rect -151 -48 -145 -14
rect -111 -48 -105 -14
rect -151 -86 -105 -48
rect -151 -120 -145 -86
rect -111 -120 -105 -86
rect -151 -158 -105 -120
rect -151 -192 -145 -158
rect -111 -192 -105 -158
rect -151 -230 -105 -192
rect -151 -264 -145 -230
rect -111 -264 -105 -230
rect -151 -302 -105 -264
rect -151 -336 -145 -302
rect -111 -336 -105 -302
rect -151 -381 -105 -336
rect -23 274 23 319
rect -23 240 -17 274
rect 17 240 23 274
rect -23 202 23 240
rect -23 168 -17 202
rect 17 168 23 202
rect -23 130 23 168
rect -23 96 -17 130
rect 17 96 23 130
rect -23 58 23 96
rect -23 24 -17 58
rect 17 24 23 58
rect -23 -14 23 24
rect -23 -48 -17 -14
rect 17 -48 23 -14
rect -23 -86 23 -48
rect -23 -120 -17 -86
rect 17 -120 23 -86
rect -23 -158 23 -120
rect -23 -192 -17 -158
rect 17 -192 23 -158
rect -23 -230 23 -192
rect -23 -264 -17 -230
rect 17 -264 23 -230
rect -23 -302 23 -264
rect -23 -336 -17 -302
rect 17 -336 23 -302
rect -23 -381 23 -336
rect 105 274 151 319
rect 105 240 111 274
rect 145 240 151 274
rect 105 202 151 240
rect 105 168 111 202
rect 145 168 151 202
rect 105 130 151 168
rect 105 96 111 130
rect 145 96 151 130
rect 105 58 151 96
rect 105 24 111 58
rect 145 24 151 58
rect 105 -14 151 24
rect 105 -48 111 -14
rect 145 -48 151 -14
rect 105 -86 151 -48
rect 105 -120 111 -86
rect 145 -120 151 -86
rect 105 -158 151 -120
rect 105 -192 111 -158
rect 145 -192 151 -158
rect 105 -230 151 -192
rect 105 -264 111 -230
rect 145 -264 151 -230
rect 105 -302 151 -264
rect 105 -336 111 -302
rect 145 -336 151 -302
rect 105 -381 151 -336
rect 233 274 279 319
rect 233 240 239 274
rect 273 240 279 274
rect 233 202 279 240
rect 233 168 239 202
rect 273 168 279 202
rect 233 130 279 168
rect 233 96 239 130
rect 273 96 279 130
rect 233 58 279 96
rect 233 24 239 58
rect 273 24 279 58
rect 233 -14 279 24
rect 233 -48 239 -14
rect 273 -48 279 -14
rect 233 -86 279 -48
rect 233 -120 239 -86
rect 273 -120 279 -86
rect 233 -158 279 -120
rect 233 -192 239 -158
rect 273 -192 279 -158
rect 233 -230 279 -192
rect 233 -264 239 -230
rect 273 -264 279 -230
rect 233 -302 279 -264
rect 233 -336 239 -302
rect 273 -336 279 -302
rect 233 -381 279 -336
rect 361 274 407 319
rect 361 240 367 274
rect 401 240 407 274
rect 361 202 407 240
rect 361 168 367 202
rect 401 168 407 202
rect 361 130 407 168
rect 361 96 367 130
rect 401 96 407 130
rect 361 58 407 96
rect 361 24 367 58
rect 401 24 407 58
rect 361 -14 407 24
rect 361 -48 367 -14
rect 401 -48 407 -14
rect 361 -86 407 -48
rect 361 -120 367 -86
rect 401 -120 407 -86
rect 361 -158 407 -120
rect 361 -192 367 -158
rect 401 -192 407 -158
rect 361 -230 407 -192
rect 361 -264 367 -230
rect 401 -264 407 -230
rect 361 -302 407 -264
rect 361 -336 367 -302
rect 401 -336 407 -302
rect 361 -381 407 -336
rect 489 274 535 319
rect 489 240 495 274
rect 529 240 535 274
rect 489 202 535 240
rect 489 168 495 202
rect 529 168 535 202
rect 489 130 535 168
rect 489 96 495 130
rect 529 96 535 130
rect 489 58 535 96
rect 489 24 495 58
rect 529 24 535 58
rect 489 -14 535 24
rect 489 -48 495 -14
rect 529 -48 535 -14
rect 489 -86 535 -48
rect 489 -120 495 -86
rect 529 -120 535 -86
rect 489 -158 535 -120
rect 489 -192 495 -158
rect 529 -192 535 -158
rect 489 -230 535 -192
rect 489 -264 495 -230
rect 529 -264 535 -230
rect 489 -302 535 -264
rect 489 -336 495 -302
rect 529 -336 535 -302
rect 489 -381 535 -336
rect 617 274 663 319
rect 617 240 623 274
rect 657 240 663 274
rect 617 202 663 240
rect 617 168 623 202
rect 657 168 663 202
rect 617 130 663 168
rect 617 96 623 130
rect 657 96 663 130
rect 617 58 663 96
rect 617 24 623 58
rect 657 24 663 58
rect 617 -14 663 24
rect 617 -48 623 -14
rect 657 -48 663 -14
rect 617 -86 663 -48
rect 617 -120 623 -86
rect 657 -120 663 -86
rect 617 -158 663 -120
rect 617 -192 623 -158
rect 657 -192 663 -158
rect 617 -230 663 -192
rect 617 -264 623 -230
rect 657 -264 663 -230
rect 617 -302 663 -264
rect 617 -336 623 -302
rect 657 -336 663 -302
rect 617 -381 663 -336
rect 745 274 791 319
rect 745 240 751 274
rect 785 240 791 274
rect 745 202 791 240
rect 745 168 751 202
rect 785 168 791 202
rect 745 130 791 168
rect 745 96 751 130
rect 785 96 791 130
rect 745 58 791 96
rect 745 24 751 58
rect 785 24 791 58
rect 745 -14 791 24
rect 745 -48 751 -14
rect 785 -48 791 -14
rect 745 -86 791 -48
rect 745 -120 751 -86
rect 785 -120 791 -86
rect 745 -158 791 -120
rect 745 -192 751 -158
rect 785 -192 791 -158
rect 745 -230 791 -192
rect 745 -264 751 -230
rect 785 -264 791 -230
rect 745 -302 791 -264
rect 745 -336 751 -302
rect 785 -336 791 -302
rect 745 -381 791 -336
rect 873 274 919 319
rect 873 240 879 274
rect 913 240 919 274
rect 873 202 919 240
rect 873 168 879 202
rect 913 168 919 202
rect 873 130 919 168
rect 873 96 879 130
rect 913 96 919 130
rect 873 58 919 96
rect 873 24 879 58
rect 913 24 919 58
rect 873 -14 919 24
rect 873 -48 879 -14
rect 913 -48 919 -14
rect 873 -86 919 -48
rect 873 -120 879 -86
rect 913 -120 919 -86
rect 873 -158 919 -120
rect 873 -192 879 -158
rect 913 -192 919 -158
rect 873 -230 919 -192
rect 873 -264 879 -230
rect 913 -264 919 -230
rect 873 -302 919 -264
rect 873 -336 879 -302
rect 913 -336 919 -302
rect 873 -381 919 -336
rect 1001 274 1047 319
rect 1001 240 1007 274
rect 1041 240 1047 274
rect 1001 202 1047 240
rect 1001 168 1007 202
rect 1041 168 1047 202
rect 1001 130 1047 168
rect 1001 96 1007 130
rect 1041 96 1047 130
rect 1001 58 1047 96
rect 1001 24 1007 58
rect 1041 24 1047 58
rect 1001 -14 1047 24
rect 1001 -48 1007 -14
rect 1041 -48 1047 -14
rect 1001 -86 1047 -48
rect 1001 -120 1007 -86
rect 1041 -120 1047 -86
rect 1001 -158 1047 -120
rect 1001 -192 1007 -158
rect 1041 -192 1047 -158
rect 1001 -230 1047 -192
rect 1001 -264 1007 -230
rect 1041 -264 1047 -230
rect 1001 -302 1047 -264
rect 1001 -336 1007 -302
rect 1041 -336 1047 -302
rect 1001 -381 1047 -336
rect 1129 274 1175 319
rect 1129 240 1135 274
rect 1169 240 1175 274
rect 1129 202 1175 240
rect 1129 168 1135 202
rect 1169 168 1175 202
rect 1129 130 1175 168
rect 1129 96 1135 130
rect 1169 96 1175 130
rect 1129 58 1175 96
rect 1129 24 1135 58
rect 1169 24 1175 58
rect 1129 -14 1175 24
rect 1129 -48 1135 -14
rect 1169 -48 1175 -14
rect 1129 -86 1175 -48
rect 1129 -120 1135 -86
rect 1169 -120 1175 -86
rect 1129 -158 1175 -120
rect 1129 -192 1135 -158
rect 1169 -192 1175 -158
rect 1129 -230 1175 -192
rect 1129 -264 1135 -230
rect 1169 -264 1175 -230
rect 1129 -302 1175 -264
rect 1129 -336 1135 -302
rect 1169 -336 1175 -302
rect 1129 -381 1175 -336
rect 1257 274 1303 319
rect 1257 240 1263 274
rect 1297 240 1303 274
rect 1257 202 1303 240
rect 1257 168 1263 202
rect 1297 168 1303 202
rect 1257 130 1303 168
rect 1257 96 1263 130
rect 1297 96 1303 130
rect 1257 58 1303 96
rect 1257 24 1263 58
rect 1297 24 1303 58
rect 1257 -14 1303 24
rect 1257 -48 1263 -14
rect 1297 -48 1303 -14
rect 1257 -86 1303 -48
rect 1257 -120 1263 -86
rect 1297 -120 1303 -86
rect 1257 -158 1303 -120
rect 1257 -192 1263 -158
rect 1297 -192 1303 -158
rect 1257 -230 1303 -192
rect 1257 -264 1263 -230
rect 1297 -264 1303 -230
rect 1257 -302 1303 -264
rect 1257 -336 1263 -302
rect 1297 -336 1303 -302
rect 1257 -381 1303 -336
rect 1385 274 1431 319
rect 1385 240 1391 274
rect 1425 240 1431 274
rect 1385 202 1431 240
rect 1385 168 1391 202
rect 1425 168 1431 202
rect 1385 130 1431 168
rect 1385 96 1391 130
rect 1425 96 1431 130
rect 1385 58 1431 96
rect 1385 24 1391 58
rect 1425 24 1431 58
rect 1385 -14 1431 24
rect 1385 -48 1391 -14
rect 1425 -48 1431 -14
rect 1385 -86 1431 -48
rect 1385 -120 1391 -86
rect 1425 -120 1431 -86
rect 1385 -158 1431 -120
rect 1385 -192 1391 -158
rect 1425 -192 1431 -158
rect 1385 -230 1431 -192
rect 1385 -264 1391 -230
rect 1425 -264 1431 -230
rect 1385 -302 1431 -264
rect 1385 -336 1391 -302
rect 1425 -336 1431 -302
rect 1385 -381 1431 -336
rect 1513 274 1559 319
rect 1513 240 1519 274
rect 1553 240 1559 274
rect 1513 202 1559 240
rect 1513 168 1519 202
rect 1553 168 1559 202
rect 1513 130 1559 168
rect 1513 96 1519 130
rect 1553 96 1559 130
rect 1513 58 1559 96
rect 1513 24 1519 58
rect 1553 24 1559 58
rect 1513 -14 1559 24
rect 1513 -48 1519 -14
rect 1553 -48 1559 -14
rect 1513 -86 1559 -48
rect 1513 -120 1519 -86
rect 1553 -120 1559 -86
rect 1513 -158 1559 -120
rect 1513 -192 1519 -158
rect 1553 -192 1559 -158
rect 1513 -230 1559 -192
rect 1513 -264 1519 -230
rect 1553 -264 1559 -230
rect 1513 -302 1559 -264
rect 1513 -336 1519 -302
rect 1553 -336 1559 -302
rect 1513 -381 1559 -336
rect 1641 274 1687 319
rect 1641 240 1647 274
rect 1681 240 1687 274
rect 1641 202 1687 240
rect 1641 168 1647 202
rect 1681 168 1687 202
rect 1641 130 1687 168
rect 1641 96 1647 130
rect 1681 96 1687 130
rect 1641 58 1687 96
rect 1641 24 1647 58
rect 1681 24 1687 58
rect 1641 -14 1687 24
rect 1641 -48 1647 -14
rect 1681 -48 1687 -14
rect 1641 -86 1687 -48
rect 1641 -120 1647 -86
rect 1681 -120 1687 -86
rect 1641 -158 1687 -120
rect 1641 -192 1647 -158
rect 1681 -192 1687 -158
rect 1641 -230 1687 -192
rect 1641 -264 1647 -230
rect 1681 -264 1687 -230
rect 1641 -302 1687 -264
rect 1641 -336 1647 -302
rect 1681 -336 1687 -302
rect 1641 -381 1687 -336
rect 1769 274 1815 319
rect 1769 240 1775 274
rect 1809 240 1815 274
rect 1769 202 1815 240
rect 1769 168 1775 202
rect 1809 168 1815 202
rect 1769 130 1815 168
rect 1769 96 1775 130
rect 1809 96 1815 130
rect 1769 58 1815 96
rect 1769 24 1775 58
rect 1809 24 1815 58
rect 1769 -14 1815 24
rect 1769 -48 1775 -14
rect 1809 -48 1815 -14
rect 1769 -86 1815 -48
rect 1769 -120 1775 -86
rect 1809 -120 1815 -86
rect 1769 -158 1815 -120
rect 1769 -192 1775 -158
rect 1809 -192 1815 -158
rect 1769 -230 1815 -192
rect 1769 -264 1775 -230
rect 1809 -264 1815 -230
rect 1769 -302 1815 -264
rect 1769 -336 1775 -302
rect 1809 -336 1815 -302
rect 1769 -381 1815 -336
rect 1897 274 1943 319
rect 1897 240 1903 274
rect 1937 240 1943 274
rect 1897 202 1943 240
rect 1897 168 1903 202
rect 1937 168 1943 202
rect 1897 130 1943 168
rect 1897 96 1903 130
rect 1937 96 1943 130
rect 1897 58 1943 96
rect 1897 24 1903 58
rect 1937 24 1943 58
rect 1897 -14 1943 24
rect 1897 -48 1903 -14
rect 1937 -48 1943 -14
rect 1897 -86 1943 -48
rect 1897 -120 1903 -86
rect 1937 -120 1943 -86
rect 1897 -158 1943 -120
rect 1897 -192 1903 -158
rect 1937 -192 1943 -158
rect 1897 -230 1943 -192
rect 1897 -264 1903 -230
rect 1937 -264 1943 -230
rect 1897 -302 1943 -264
rect 1897 -336 1903 -302
rect 1937 -336 1943 -302
rect 1897 -381 1943 -336
rect 2025 274 2071 319
rect 2025 240 2031 274
rect 2065 240 2071 274
rect 2025 202 2071 240
rect 2025 168 2031 202
rect 2065 168 2071 202
rect 2025 130 2071 168
rect 2025 96 2031 130
rect 2065 96 2071 130
rect 2025 58 2071 96
rect 2025 24 2031 58
rect 2065 24 2071 58
rect 2025 -14 2071 24
rect 2025 -48 2031 -14
rect 2065 -48 2071 -14
rect 2025 -86 2071 -48
rect 2025 -120 2031 -86
rect 2065 -120 2071 -86
rect 2025 -158 2071 -120
rect 2025 -192 2031 -158
rect 2065 -192 2071 -158
rect 2025 -230 2071 -192
rect 2025 -264 2031 -230
rect 2065 -264 2071 -230
rect 2025 -302 2071 -264
rect 2025 -336 2031 -302
rect 2065 -336 2071 -302
rect 2025 -381 2071 -336
<< labels >>
flabel metal1 s -1984 374 -1984 374 0 FreeSans 300 0 0 0 G
port 1 nsew
flabel metal1 s -1855 374 -1855 374 0 FreeSans 300 0 0 0 G
port 1 nsew
flabel metal1 s -1728 374 -1728 374 0 FreeSans 300 0 0 0 G
port 1 nsew
flabel metal1 s -1600 374 -1600 374 0 FreeSans 300 0 0 0 G
port 1 nsew
flabel metal1 s -1472 374 -1472 374 0 FreeSans 300 0 0 0 G
port 1 nsew
flabel metal1 s -1344 374 -1344 374 0 FreeSans 300 0 0 0 G
port 1 nsew
flabel metal1 s -1216 374 -1216 374 0 FreeSans 300 0 0 0 G
port 1 nsew
flabel metal1 s -1088 374 -1088 374 0 FreeSans 300 0 0 0 G
port 1 nsew
flabel metal1 s -960 374 -960 374 0 FreeSans 300 0 0 0 G
port 1 nsew
flabel metal1 s -832 374 -832 374 0 FreeSans 300 0 0 0 G
port 1 nsew
flabel metal1 s -704 374 -704 374 0 FreeSans 300 0 0 0 G
port 1 nsew
flabel metal1 s -576 374 -576 374 0 FreeSans 300 0 0 0 G
port 1 nsew
flabel metal1 s -448 374 -448 374 0 FreeSans 300 0 0 0 G
port 1 nsew
flabel metal1 s -320 374 -320 374 0 FreeSans 300 0 0 0 G
port 1 nsew
flabel metal1 s -192 374 -192 374 0 FreeSans 300 0 0 0 G
port 1 nsew
flabel metal1 s -64 374 -64 374 0 FreeSans 300 0 0 0 G
port 1 nsew
flabel metal1 s 64 374 64 374 0 FreeSans 300 0 0 0 G
port 1 nsew
flabel metal1 s 192 374 192 374 0 FreeSans 300 0 0 0 G
port 1 nsew
flabel metal1 s 320 374 320 374 0 FreeSans 300 0 0 0 G
port 1 nsew
flabel metal1 s 448 374 448 374 0 FreeSans 300 0 0 0 G
port 1 nsew
flabel metal1 s 576 374 576 374 0 FreeSans 300 0 0 0 G
port 1 nsew
flabel metal1 s 704 374 704 374 0 FreeSans 300 0 0 0 G
port 1 nsew
flabel metal1 s 832 374 832 374 0 FreeSans 300 0 0 0 G
port 1 nsew
flabel metal1 s 960 374 960 374 0 FreeSans 300 0 0 0 G
port 1 nsew
flabel metal1 s 1088 374 1088 374 0 FreeSans 300 0 0 0 G
port 1 nsew
flabel metal1 s 1216 374 1216 374 0 FreeSans 300 0 0 0 G
port 1 nsew
flabel metal1 s 1344 374 1344 374 0 FreeSans 300 0 0 0 G
port 1 nsew
flabel metal1 s 1472 374 1472 374 0 FreeSans 300 0 0 0 G
port 1 nsew
flabel metal1 s 1600 374 1600 374 0 FreeSans 300 0 0 0 G
port 1 nsew
flabel metal1 s 1728 374 1728 374 0 FreeSans 300 0 0 0 G
port 1 nsew
flabel metal1 s 1855 374 1855 374 0 FreeSans 300 0 0 0 G
port 1 nsew
flabel metal1 s 1984 374 1984 374 0 FreeSans 300 0 0 0 G
port 1 nsew
flabel metal1 s -2048 -31 -2048 -31 0 FreeSans 300 0 0 0 D
port 2 nsew
flabel metal1 s -1920 -31 -1920 -31 0 FreeSans 300 0 0 0 S
port 3 nsew
flabel metal1 s -1792 -31 -1792 -31 0 FreeSans 300 0 0 0 D
port 2 nsew
flabel metal1 s -1664 -31 -1664 -31 0 FreeSans 300 0 0 0 S
port 3 nsew
flabel metal1 s -1536 -31 -1536 -31 0 FreeSans 300 0 0 0 D
port 2 nsew
flabel metal1 s -1408 -31 -1408 -31 0 FreeSans 300 0 0 0 S
port 3 nsew
flabel metal1 s -1280 -31 -1280 -31 0 FreeSans 300 0 0 0 D
port 2 nsew
flabel metal1 s -1152 -31 -1152 -31 0 FreeSans 300 0 0 0 S
port 3 nsew
flabel metal1 s -1024 -31 -1024 -31 0 FreeSans 300 0 0 0 D
port 2 nsew
flabel metal1 s -896 -31 -896 -31 0 FreeSans 300 0 0 0 S
port 3 nsew
flabel metal1 s -768 -31 -768 -31 0 FreeSans 300 0 0 0 D
port 2 nsew
flabel metal1 s -640 -31 -640 -31 0 FreeSans 300 0 0 0 S
port 3 nsew
flabel metal1 s -512 -31 -512 -31 0 FreeSans 300 0 0 0 D
port 2 nsew
flabel metal1 s -384 -31 -384 -31 0 FreeSans 300 0 0 0 S
port 3 nsew
flabel metal1 s -256 -31 -256 -31 0 FreeSans 300 0 0 0 D
port 2 nsew
flabel metal1 s -128 -31 -128 -31 0 FreeSans 300 0 0 0 S
port 3 nsew
flabel metal1 s 0 -31 0 -31 0 FreeSans 300 0 0 0 D
port 2 nsew
flabel metal1 s 128 -31 128 -31 0 FreeSans 300 0 0 0 S
port 3 nsew
flabel metal1 s 256 -31 256 -31 0 FreeSans 300 0 0 0 D
port 2 nsew
flabel metal1 s 384 -31 384 -31 0 FreeSans 300 0 0 0 S
port 3 nsew
flabel metal1 s 512 -31 512 -31 0 FreeSans 300 0 0 0 D
port 2 nsew
flabel metal1 s 640 -31 640 -31 0 FreeSans 300 0 0 0 S
port 3 nsew
flabel metal1 s 768 -31 768 -31 0 FreeSans 300 0 0 0 D
port 2 nsew
flabel metal1 s 896 -31 896 -31 0 FreeSans 300 0 0 0 S
port 3 nsew
flabel metal1 s 1024 -31 1024 -31 0 FreeSans 300 0 0 0 D
port 2 nsew
flabel metal1 s 1152 -31 1152 -31 0 FreeSans 300 0 0 0 S
port 3 nsew
flabel metal1 s 1280 -31 1280 -31 0 FreeSans 300 0 0 0 D
port 2 nsew
flabel metal1 s 1408 -31 1408 -31 0 FreeSans 300 0 0 0 S
port 3 nsew
flabel metal1 s 1536 -31 1536 -31 0 FreeSans 300 0 0 0 D
port 2 nsew
flabel metal1 s 1664 -31 1664 -31 0 FreeSans 300 0 0 0 S
port 3 nsew
flabel metal1 s 1792 -31 1792 -31 0 FreeSans 300 0 0 0 D
port 2 nsew
flabel metal1 s 1920 -31 1920 -31 0 FreeSans 300 0 0 0 S
port 3 nsew
flabel metal1 s 2048 -31 2048 -31 0 FreeSans 300 0 0 0 D
port 2 nsew
<< properties >>
string FIXED_BBOX -2162 -476 2162 476
<< end >>
