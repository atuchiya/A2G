magic
tech sky130A
timestamp 1680007175
<< error_p >>
rect -5 5 5 9
rect -5 -5 9 5
<< metal1 >>
rect -5 -5 5 5
<< labels >>
<< end >>
