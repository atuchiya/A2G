magic
tech sky130A
magscale 1 2
timestamp 1686266348
<< checkpaint >>
rect -1899 -1624 1899 1624
<< nwell >>
rect -639 -364 639 364
<< pmos >>
rect -443 -216 -383 144
rect -325 -216 -265 144
rect -207 -216 -147 144
rect -89 -216 -29 144
rect 29 -216 89 144
rect 147 -216 207 144
rect 265 -216 325 144
rect 383 -216 443 144
<< pdiff >>
rect -501 132 -443 144
rect -501 -204 -489 132
rect -455 -204 -443 132
rect -501 -216 -443 -204
rect -383 132 -325 144
rect -383 -204 -371 132
rect -337 -204 -325 132
rect -383 -216 -325 -204
rect -265 132 -207 144
rect -265 -204 -253 132
rect -219 -204 -207 132
rect -265 -216 -207 -204
rect -147 132 -89 144
rect -147 -204 -135 132
rect -101 -204 -89 132
rect -147 -216 -89 -204
rect -29 132 29 144
rect -29 -204 -17 132
rect 17 -204 29 132
rect -29 -216 29 -204
rect 89 132 147 144
rect 89 -204 101 132
rect 135 -204 147 132
rect 89 -216 147 -204
rect 207 132 265 144
rect 207 -204 219 132
rect 253 -204 265 132
rect 207 -216 265 -204
rect 325 132 383 144
rect 325 -204 337 132
rect 371 -204 383 132
rect 325 -216 383 -204
rect 443 132 501 144
rect 443 -204 455 132
rect 489 -204 501 132
rect 443 -216 501 -204
<< pdiffc >>
rect -489 -204 -455 132
rect -371 -204 -337 132
rect -253 -204 -219 132
rect -135 -204 -101 132
rect -17 -204 17 132
rect 101 -204 135 132
rect 219 -204 253 132
rect 337 -204 371 132
rect 455 -204 489 132
<< nsubdiff >>
rect -603 294 -507 328
rect 507 294 603 328
rect -603 231 -569 294
rect 569 231 603 294
rect -603 -294 -569 -231
rect 569 -294 603 -231
rect -603 -328 -507 -294
rect 507 -328 603 -294
<< nsubdiffcont >>
rect -507 294 507 328
rect -603 -231 -569 231
rect 569 -231 603 231
rect -507 -328 507 -294
<< poly >>
rect -446 225 -380 241
rect -446 191 -430 225
rect -396 191 -380 225
rect -446 175 -380 191
rect -328 225 -262 241
rect -328 191 -312 225
rect -278 191 -262 225
rect -328 175 -262 191
rect -210 225 -144 241
rect -210 191 -194 225
rect -160 191 -144 225
rect -210 175 -144 191
rect -92 225 -26 241
rect -92 191 -76 225
rect -42 191 -26 225
rect -92 175 -26 191
rect 26 225 92 241
rect 26 191 42 225
rect 76 191 92 225
rect 26 175 92 191
rect 144 225 210 241
rect 144 191 160 225
rect 194 191 210 225
rect 144 175 210 191
rect 262 225 328 241
rect 262 191 278 225
rect 312 191 328 225
rect 262 175 328 191
rect 380 225 446 241
rect 380 191 396 225
rect 430 191 446 225
rect 380 175 446 191
rect -443 144 -383 175
rect -325 144 -265 175
rect -207 144 -147 175
rect -89 144 -29 175
rect 29 144 89 175
rect 147 144 207 175
rect 265 144 325 175
rect 383 144 443 175
rect -443 -242 -383 -216
rect -325 -242 -265 -216
rect -207 -242 -147 -216
rect -89 -242 -29 -216
rect 29 -242 89 -216
rect 147 -242 207 -216
rect 265 -242 325 -216
rect 383 -242 443 -216
<< polycont >>
rect -430 191 -396 225
rect -312 191 -278 225
rect -194 191 -160 225
rect -76 191 -42 225
rect 42 191 76 225
rect 160 191 194 225
rect 278 191 312 225
rect 396 191 430 225
<< locali >>
rect -603 294 -507 328
rect 507 294 603 328
rect -603 231 -569 294
rect 569 231 603 294
rect -446 191 -430 225
rect -396 191 -380 225
rect -328 191 -312 225
rect -278 191 -262 225
rect -210 191 -194 225
rect -160 191 -144 225
rect -92 191 -76 225
rect -42 191 -26 225
rect 26 191 42 225
rect 76 191 92 225
rect 144 191 160 225
rect 194 191 210 225
rect 262 191 278 225
rect 312 191 328 225
rect 380 191 396 225
rect 430 191 446 225
rect -489 132 -455 148
rect -489 -220 -455 -204
rect -371 132 -337 148
rect -371 -220 -337 -204
rect -253 132 -219 148
rect -253 -220 -219 -204
rect -135 132 -101 148
rect -135 -220 -101 -204
rect -17 132 17 148
rect -17 -220 17 -204
rect 101 132 135 148
rect 101 -220 135 -204
rect 219 132 253 148
rect 219 -220 253 -204
rect 337 132 371 148
rect 337 -220 371 -204
rect 455 132 489 148
rect 455 -220 489 -204
rect -603 -294 -569 -231
rect 569 -294 603 -231
rect -603 -328 -507 -294
rect 507 -328 603 -294
<< viali >>
rect -430 191 -396 225
rect -312 191 -278 225
rect -194 191 -160 225
rect -76 191 -42 225
rect 42 191 76 225
rect 160 191 194 225
rect 278 191 312 225
rect 396 191 430 225
rect -489 -204 -455 132
rect -371 -204 -337 132
rect -253 -204 -219 132
rect -135 -204 -101 132
rect -17 -204 17 132
rect 101 -204 135 132
rect 219 -204 253 132
rect 337 -204 371 132
rect 455 -204 489 132
<< metal1 >>
rect -442 225 -384 231
rect -442 191 -430 225
rect -396 191 -384 225
rect -442 185 -384 191
rect -324 225 -266 231
rect -324 191 -312 225
rect -278 191 -266 225
rect -324 185 -266 191
rect -206 225 -148 231
rect -206 191 -194 225
rect -160 191 -148 225
rect -206 185 -148 191
rect -88 225 -30 231
rect -88 191 -76 225
rect -42 191 -30 225
rect -88 185 -30 191
rect 30 225 88 231
rect 30 191 42 225
rect 76 191 88 225
rect 30 185 88 191
rect 148 225 206 231
rect 148 191 160 225
rect 194 191 206 225
rect 148 185 206 191
rect 266 225 324 231
rect 266 191 278 225
rect 312 191 324 225
rect 266 185 324 191
rect 384 225 442 231
rect 384 191 396 225
rect 430 191 442 225
rect 384 185 442 191
rect -495 132 -449 144
rect -495 -204 -489 132
rect -455 -204 -449 132
rect -495 -216 -449 -204
rect -377 132 -331 144
rect -377 -204 -371 132
rect -337 -204 -331 132
rect -377 -216 -331 -204
rect -259 132 -213 144
rect -259 -204 -253 132
rect -219 -204 -213 132
rect -259 -216 -213 -204
rect -141 132 -95 144
rect -141 -204 -135 132
rect -101 -204 -95 132
rect -141 -216 -95 -204
rect -23 132 23 144
rect -23 -204 -17 132
rect 17 -204 23 132
rect -23 -216 23 -204
rect 95 132 141 144
rect 95 -204 101 132
rect 135 -204 141 132
rect 95 -216 141 -204
rect 213 132 259 144
rect 213 -204 219 132
rect 253 -204 259 132
rect 213 -216 259 -204
rect 331 132 377 144
rect 331 -204 337 132
rect 371 -204 377 132
rect 331 -216 377 -204
rect 449 132 495 144
rect 449 -204 455 132
rect 489 -204 495 132
rect 449 -216 495 -204
<< labels >>
flabel metal1 -413 208 -413 208 0 FreeSans 240 0 0 0 G
flabel metal1 -295 208 -295 208 0 FreeSans 240 0 0 0 G
flabel metal1 -177 208 -177 208 0 FreeSans 240 0 0 0 G
flabel metal1 -59 208 -59 208 0 FreeSans 240 0 0 0 G
flabel metal1 59 208 59 208 0 FreeSans 240 0 0 0 G
flabel metal1 177 208 177 208 0 FreeSans 240 0 0 0 G
flabel metal1 295 208 295 208 0 FreeSans 240 0 0 0 G
flabel metal1 413 208 413 208 0 FreeSans 240 0 0 0 G
flabel metal1 -472 -36 -472 -36 0 FreeSans 240 0 0 0 D
flabel metal1 -354 -36 -354 -36 0 FreeSans 240 0 0 0 S
flabel metal1 -236 -36 -236 -36 0 FreeSans 240 0 0 0 D
flabel metal1 -118 -36 -118 -36 0 FreeSans 240 0 0 0 S
flabel metal1 0 -36 0 -36 0 FreeSans 240 0 0 0 D
flabel metal1 118 -36 118 -36 0 FreeSans 240 0 0 0 S
flabel metal1 236 -36 236 -36 0 FreeSans 240 0 0 0 D
flabel metal1 354 -36 354 -36 0 FreeSans 240 0 0 0 S
flabel metal1 472 -36 472 -36 0 FreeSans 240 0 0 0 D
<< properties >>
string FIXED_BBOX -586 -311 586 311
<< end >>

