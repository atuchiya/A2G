magic
tech sky130A
magscale 1 2
timestamp 1686266346
<< checkpaint >>
rect -2135 -1619 2135 1619
<< pwell >>
rect -875 -359 875 359
<< nmos >>
rect -679 -211 -619 149
rect -561 -211 -501 149
rect -443 -211 -383 149
rect -325 -211 -265 149
rect -207 -211 -147 149
rect -89 -211 -29 149
rect 29 -211 89 149
rect 147 -211 207 149
rect 265 -211 325 149
rect 383 -211 443 149
rect 501 -211 561 149
rect 619 -211 679 149
<< ndiff >>
rect -737 137 -679 149
rect -737 -199 -725 137
rect -691 -199 -679 137
rect -737 -211 -679 -199
rect -619 137 -561 149
rect -619 -199 -607 137
rect -573 -199 -561 137
rect -619 -211 -561 -199
rect -501 137 -443 149
rect -501 -199 -489 137
rect -455 -199 -443 137
rect -501 -211 -443 -199
rect -383 137 -325 149
rect -383 -199 -371 137
rect -337 -199 -325 137
rect -383 -211 -325 -199
rect -265 137 -207 149
rect -265 -199 -253 137
rect -219 -199 -207 137
rect -265 -211 -207 -199
rect -147 137 -89 149
rect -147 -199 -135 137
rect -101 -199 -89 137
rect -147 -211 -89 -199
rect -29 137 29 149
rect -29 -199 -17 137
rect 17 -199 29 137
rect -29 -211 29 -199
rect 89 137 147 149
rect 89 -199 101 137
rect 135 -199 147 137
rect 89 -211 147 -199
rect 207 137 265 149
rect 207 -199 219 137
rect 253 -199 265 137
rect 207 -211 265 -199
rect 325 137 383 149
rect 325 -199 337 137
rect 371 -199 383 137
rect 325 -211 383 -199
rect 443 137 501 149
rect 443 -199 455 137
rect 489 -199 501 137
rect 443 -211 501 -199
rect 561 137 619 149
rect 561 -199 573 137
rect 607 -199 619 137
rect 561 -211 619 -199
rect 679 137 737 149
rect 679 -199 691 137
rect 725 -199 737 137
rect 679 -211 737 -199
<< ndiffc >>
rect -725 -199 -691 137
rect -607 -199 -573 137
rect -489 -199 -455 137
rect -371 -199 -337 137
rect -253 -199 -219 137
rect -135 -199 -101 137
rect -17 -199 17 137
rect 101 -199 135 137
rect 219 -199 253 137
rect 337 -199 371 137
rect 455 -199 489 137
rect 573 -199 607 137
rect 691 -199 725 137
<< psubdiff >>
rect -839 289 -743 323
rect 743 289 839 323
rect -839 227 -805 289
rect 805 227 839 289
rect -839 -289 -805 -227
rect 805 -289 839 -227
rect -839 -323 -743 -289
rect 743 -323 839 -289
<< psubdiffcont >>
rect -743 289 743 323
rect -839 -227 -805 227
rect 805 -227 839 227
rect -743 -323 743 -289
<< poly >>
rect -682 221 -616 237
rect -682 187 -666 221
rect -632 187 -616 221
rect -682 171 -616 187
rect -564 221 -498 237
rect -564 187 -548 221
rect -514 187 -498 221
rect -564 171 -498 187
rect -446 221 -380 237
rect -446 187 -430 221
rect -396 187 -380 221
rect -446 171 -380 187
rect -328 221 -262 237
rect -328 187 -312 221
rect -278 187 -262 221
rect -328 171 -262 187
rect -210 221 -144 237
rect -210 187 -194 221
rect -160 187 -144 221
rect -210 171 -144 187
rect -92 221 -26 237
rect -92 187 -76 221
rect -42 187 -26 221
rect -92 171 -26 187
rect 26 221 92 237
rect 26 187 42 221
rect 76 187 92 221
rect 26 171 92 187
rect 144 221 210 237
rect 144 187 160 221
rect 194 187 210 221
rect 144 171 210 187
rect 262 221 328 237
rect 262 187 278 221
rect 312 187 328 221
rect 262 171 328 187
rect 380 221 446 237
rect 380 187 396 221
rect 430 187 446 221
rect 380 171 446 187
rect 498 221 564 237
rect 498 187 514 221
rect 548 187 564 221
rect 498 171 564 187
rect 616 221 682 237
rect 616 187 632 221
rect 666 187 682 221
rect 616 171 682 187
rect -679 149 -619 171
rect -561 149 -501 171
rect -443 149 -383 171
rect -325 149 -265 171
rect -207 149 -147 171
rect -89 149 -29 171
rect 29 149 89 171
rect 147 149 207 171
rect 265 149 325 171
rect 383 149 443 171
rect 501 149 561 171
rect 619 149 679 171
rect -679 -237 -619 -211
rect -561 -237 -501 -211
rect -443 -237 -383 -211
rect -325 -237 -265 -211
rect -207 -237 -147 -211
rect -89 -237 -29 -211
rect 29 -237 89 -211
rect 147 -237 207 -211
rect 265 -237 325 -211
rect 383 -237 443 -211
rect 501 -237 561 -211
rect 619 -237 679 -211
<< polycont >>
rect -666 187 -632 221
rect -548 187 -514 221
rect -430 187 -396 221
rect -312 187 -278 221
rect -194 187 -160 221
rect -76 187 -42 221
rect 42 187 76 221
rect 160 187 194 221
rect 278 187 312 221
rect 396 187 430 221
rect 514 187 548 221
rect 632 187 666 221
<< locali >>
rect -839 289 -743 323
rect 743 289 839 323
rect -839 227 -805 289
rect 805 227 839 289
rect -682 187 -666 221
rect -632 187 -616 221
rect -564 187 -548 221
rect -514 187 -498 221
rect -446 187 -430 221
rect -396 187 -380 221
rect -328 187 -312 221
rect -278 187 -262 221
rect -210 187 -194 221
rect -160 187 -144 221
rect -92 187 -76 221
rect -42 187 -26 221
rect 26 187 42 221
rect 76 187 92 221
rect 144 187 160 221
rect 194 187 210 221
rect 262 187 278 221
rect 312 187 328 221
rect 380 187 396 221
rect 430 187 446 221
rect 498 187 514 221
rect 548 187 564 221
rect 616 187 632 221
rect 666 187 682 221
rect -725 137 -691 153
rect -725 -215 -691 -199
rect -607 137 -573 153
rect -607 -215 -573 -199
rect -489 137 -455 153
rect -489 -215 -455 -199
rect -371 137 -337 153
rect -371 -215 -337 -199
rect -253 137 -219 153
rect -253 -215 -219 -199
rect -135 137 -101 153
rect -135 -215 -101 -199
rect -17 137 17 153
rect -17 -215 17 -199
rect 101 137 135 153
rect 101 -215 135 -199
rect 219 137 253 153
rect 219 -215 253 -199
rect 337 137 371 153
rect 337 -215 371 -199
rect 455 137 489 153
rect 455 -215 489 -199
rect 573 137 607 153
rect 573 -215 607 -199
rect 691 137 725 153
rect 691 -215 725 -199
rect -839 -289 -805 -227
rect 805 -289 839 -227
rect -839 -323 -743 -289
rect 743 -323 839 -289
<< viali >>
rect -666 187 -632 221
rect -548 187 -514 221
rect -430 187 -396 221
rect -312 187 -278 221
rect -194 187 -160 221
rect -76 187 -42 221
rect 42 187 76 221
rect 160 187 194 221
rect 278 187 312 221
rect 396 187 430 221
rect 514 187 548 221
rect 632 187 666 221
rect -725 -199 -691 137
rect -607 -199 -573 137
rect -489 -199 -455 137
rect -371 -199 -337 137
rect -253 -199 -219 137
rect -135 -199 -101 137
rect -17 -199 17 137
rect 101 -199 135 137
rect 219 -199 253 137
rect 337 -199 371 137
rect 455 -199 489 137
rect 573 -199 607 137
rect 691 -199 725 137
<< metal1 >>
rect -678 221 -620 227
rect -678 187 -666 221
rect -632 187 -620 221
rect -678 181 -620 187
rect -560 221 -502 227
rect -560 187 -548 221
rect -514 187 -502 221
rect -560 181 -502 187
rect -442 221 -384 227
rect -442 187 -430 221
rect -396 187 -384 221
rect -442 181 -384 187
rect -324 221 -266 227
rect -324 187 -312 221
rect -278 187 -266 221
rect -324 181 -266 187
rect -206 221 -148 227
rect -206 187 -194 221
rect -160 187 -148 221
rect -206 181 -148 187
rect -88 221 -30 227
rect -88 187 -76 221
rect -42 187 -30 221
rect -88 181 -30 187
rect 30 221 88 227
rect 30 187 42 221
rect 76 187 88 221
rect 30 181 88 187
rect 148 221 206 227
rect 148 187 160 221
rect 194 187 206 221
rect 148 181 206 187
rect 266 221 324 227
rect 266 187 278 221
rect 312 187 324 221
rect 266 181 324 187
rect 384 221 442 227
rect 384 187 396 221
rect 430 187 442 221
rect 384 181 442 187
rect 502 221 560 227
rect 502 187 514 221
rect 548 187 560 221
rect 502 181 560 187
rect 620 221 678 227
rect 620 187 632 221
rect 666 187 678 221
rect 620 181 678 187
rect -731 137 -685 149
rect -731 -199 -725 137
rect -691 -199 -685 137
rect -731 -211 -685 -199
rect -613 137 -567 149
rect -613 -199 -607 137
rect -573 -199 -567 137
rect -613 -211 -567 -199
rect -495 137 -449 149
rect -495 -199 -489 137
rect -455 -199 -449 137
rect -495 -211 -449 -199
rect -377 137 -331 149
rect -377 -199 -371 137
rect -337 -199 -331 137
rect -377 -211 -331 -199
rect -259 137 -213 149
rect -259 -199 -253 137
rect -219 -199 -213 137
rect -259 -211 -213 -199
rect -141 137 -95 149
rect -141 -199 -135 137
rect -101 -199 -95 137
rect -141 -211 -95 -199
rect -23 137 23 149
rect -23 -199 -17 137
rect 17 -199 23 137
rect -23 -211 23 -199
rect 95 137 141 149
rect 95 -199 101 137
rect 135 -199 141 137
rect 95 -211 141 -199
rect 213 137 259 149
rect 213 -199 219 137
rect 253 -199 259 137
rect 213 -211 259 -199
rect 331 137 377 149
rect 331 -199 337 137
rect 371 -199 377 137
rect 331 -211 377 -199
rect 449 137 495 149
rect 449 -199 455 137
rect 489 -199 495 137
rect 449 -211 495 -199
rect 567 137 613 149
rect 567 -199 573 137
rect 607 -199 613 137
rect 567 -211 613 -199
rect 685 137 731 149
rect 685 -199 691 137
rect 725 -199 731 137
rect 685 -211 731 -199
<< labels >>
flabel metal1 -649 204 -649 204 0 FreeSans 240 0 0 0 G
flabel metal1 -531 204 -531 204 0 FreeSans 240 0 0 0 G
flabel metal1 -413 204 -413 204 0 FreeSans 240 0 0 0 G
flabel metal1 -295 204 -295 204 0 FreeSans 240 0 0 0 G
flabel metal1 -177 204 -177 204 0 FreeSans 240 0 0 0 G
flabel metal1 -59 204 -59 204 0 FreeSans 240 0 0 0 G
flabel metal1 59 204 59 204 0 FreeSans 240 0 0 0 G
flabel metal1 177 204 177 204 0 FreeSans 240 0 0 0 G
flabel metal1 295 204 295 204 0 FreeSans 240 0 0 0 G
flabel metal1 413 204 413 204 0 FreeSans 240 0 0 0 G
flabel metal1 531 204 531 204 0 FreeSans 240 0 0 0 G
flabel metal1 649 204 649 204 0 FreeSans 240 0 0 0 G
flabel metal1 -708 -31 -708 -31 0 FreeSans 240 0 0 0 D
flabel metal1 -590 -31 -590 -31 0 FreeSans 240 0 0 0 S
flabel metal1 -472 -31 -472 -31 0 FreeSans 240 0 0 0 D
flabel metal1 -354 -31 -354 -31 0 FreeSans 240 0 0 0 S
flabel metal1 -236 -31 -236 -31 0 FreeSans 240 0 0 0 D
flabel metal1 -118 -31 -118 -31 0 FreeSans 240 0 0 0 S
flabel metal1 0 -31 0 -31 0 FreeSans 240 0 0 0 D
flabel metal1 118 -31 118 -31 0 FreeSans 240 0 0 0 S
flabel metal1 236 -31 236 -31 0 FreeSans 240 0 0 0 D
flabel metal1 354 -31 354 -31 0 FreeSans 240 0 0 0 S
flabel metal1 472 -31 472 -31 0 FreeSans 240 0 0 0 D
flabel metal1 590 -31 590 -31 0 FreeSans 240 0 0 0 S
flabel metal1 708 -31 708 -31 0 FreeSans 240 0 0 0 D
<< properties >>
string FIXED_BBOX -822 -306 822 306
<< end >>

