magic
tech sky130A
magscale 1 2
timestamp 1686266350
<< checkpaint >>
rect -1899 -1619 1899 1619
<< metal2 >>
rect -444 180 444 244
rect -504 -32 504 32
rect -386 -232 386 -168
use via_M1_M2_1  NoName_177 ~/A2G/A2G/magic/magic_layout/skywater130_microtemplates_dense
timestamp 1647525606
transform 1 0 -472 0 1 0
box -32 -32 32 32
use via_M1_M2_1  NoName_178
timestamp 1647525606
transform 1 0 -236 0 1 0
box -32 -32 32 32
use via_M1_M2_1  NoName_179
timestamp 1647525606
transform 1 0 0 0 1 0
box -32 -32 32 32
use via_M1_M2_1  NoName_180
timestamp 1647525606
transform 1 0 236 0 1 0
box -32 -32 32 32
use via_M1_M2_1  NoName_181
timestamp 1647525606
transform 1 0 472 0 1 0
box -32 -32 32 32
use via_M1_M2_1  NoName_182
timestamp 1647525606
transform 1 0 -354 0 1 -200
box -32 -32 32 32
use via_M1_M2_1  NoName_183
timestamp 1647525606
transform 1 0 -118 0 1 -200
box -32 -32 32 32
use via_M1_M2_1  NoName_184
timestamp 1647525606
transform 1 0 118 0 1 -200
box -32 -32 32 32
use via_M1_M2_1  NoName_185
timestamp 1647525606
transform 1 0 354 0 1 -200
box -32 -32 32 32
use via_M1_M2_1  NoName_186
timestamp 1647525606
transform 1 0 -412 0 1 212
box -32 -32 32 32
use via_M1_M2_1  NoName_187
timestamp 1647525606
transform 1 0 -294 0 1 212
box -32 -32 32 32
use via_M1_M2_1  NoName_188
timestamp 1647525606
transform 1 0 -176 0 1 212
box -32 -32 32 32
use via_M1_M2_1  NoName_189
timestamp 1647525606
transform 1 0 -58 0 1 212
box -32 -32 32 32
use via_M1_M2_1  NoName_190
timestamp 1647525606
transform 1 0 58 0 1 212
box -32 -32 32 32
use via_M1_M2_1  NoName_191
timestamp 1647525606
transform 1 0 176 0 1 212
box -32 -32 32 32
use via_M1_M2_1  NoName_192
timestamp 1647525606
transform 1 0 294 0 1 212
box -32 -32 32 32
use via_M1_M2_1  NoName_193
timestamp 1647525606
transform 1 0 412 0 1 212
box -32 -32 32 32
use XMl2_origin  XMl2
timestamp 1686266350
transform 1 0 0 0 1 0
box -639 -359 639 359
<< end >>
