.subckt diff2sin vdd vss out ib ia icmbias
*.iopin vdd
*.iopin vss
*.opin out
*.ipin ib
*.ipin ia
*.ipin icmbias
XM1 net1 ia net2 vss sky130_fd_pr__nfet_01v8_lvt L=l W=w nf=1 ad='int((nf+1)/2) * W/nf * 0.29' as='int((nf+2)/2) * W/nf * 0.29'
+ pd='2*int((nf+1)/2) * (W/nf + 0.29)' ps='2*int((nf+2)/2) * (W/nf + 0.29)' nrd='0.29 / W' nrs='0.29 / W'
+ sa=0 sb=0 sd=0 mult=m1 m=m1
XM2 net1 net1 vdd vdd sky130_fd_pr__pfet_01v8_lvt L=l W=w nf=1 ad='int((nf+1)/2) * W/nf * 0.29' as='int((nf+2)/2) * W/nf * 0.29'
+ pd='2*int((nf+1)/2) * (W/nf + 0.29)' ps='2*int((nf+2)/2) * (W/nf + 0.29)' nrd='0.29 / W' nrs='0.29 / W'
+ sa=0 sb=0 sd=0 mult=m2 m=m2
XM3 out ib net2 vss sky130_fd_pr__nfet_01v8_lvt L=l W=w nf=1 ad='int((nf+1)/2) * W/nf * 0.29' as='int((nf+2)/2) * W/nf * 0.29'
+ pd='2*int((nf+1)/2) * (W/nf + 0.29)' ps='2*int((nf+2)/2) * (W/nf + 0.29)' nrd='0.29 / W' nrs='0.29 / W'
+ sa=0 sb=0 sd=0 mult=m3 m=m3
XM4 out net1 vdd vdd sky130_fd_pr__pfet_01v8_lvt L=l W=w nf=1 ad='int((nf+1)/2) * W/nf * 0.29' as='int((nf+2)/2) * W/nf * 0.29'
+ pd='2*int((nf+1)/2) * (W/nf + 0.29)' ps='2*int((nf+2)/2) * (W/nf + 0.29)' nrd='0.29 / W' nrs='0.29 / W'
+ sa=0 sb=0 sd=0 mult=m4 m=m4
XM5 net2 icmbias vss vss sky130_fd_pr__nfet_01v8_lvt L=l W=w nf=1 ad='int((nf+1)/2) * W/nf * 0.29' as='int((nf+2)/2) * W/nf * 0.29'
+ pd='2*int((nf+1)/2) * (W/nf + 0.29)' ps='2*int((nf+2)/2) * (W/nf + 0.29)' nrd='0.29 / W' nrs='0.29 / W'
+ sa=0 sb=0 sd=0 mult=m5 m=m5
.param w=3.5
.param l=0.35
.param m1=16
.param m2=40
.param m3=16
.param m4=40
.param m5=32
.ends
*.end