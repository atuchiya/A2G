magic
tech sky130A
magscale 1 2
timestamp 1686232357
<< checkpaint >>
rect -3987 -1794 3987 1794
<< metal2 >>
rect -2528 380 2528 444
rect -2592 -32 2592 32
rect -2464 -432 2464 -368
use via_M1_M2_1  NoName_148 ~/A2G/A2G/magic/magic_layout/skywater130_microtemplates_dense
timestamp 1647525606
transform 1 0 -2560 0 1 0
box -32 -32 32 32
use via_M1_M2_1  NoName_149
timestamp 1647525606
transform 1 0 -2304 0 1 0
box -32 -32 32 32
use via_M1_M2_1  NoName_150
timestamp 1647525606
transform 1 0 -2048 0 1 0
box -32 -32 32 32
use via_M1_M2_1  NoName_151
timestamp 1647525606
transform 1 0 -1792 0 1 0
box -32 -32 32 32
use via_M1_M2_1  NoName_152
timestamp 1647525606
transform 1 0 -1536 0 1 0
box -32 -32 32 32
use via_M1_M2_1  NoName_153
timestamp 1647525606
transform 1 0 -1280 0 1 0
box -32 -32 32 32
use via_M1_M2_1  NoName_154
timestamp 1647525606
transform 1 0 -1024 0 1 0
box -32 -32 32 32
use via_M1_M2_1  NoName_155
timestamp 1647525606
transform 1 0 -768 0 1 0
box -32 -32 32 32
use via_M1_M2_1  NoName_156
timestamp 1647525606
transform 1 0 -512 0 1 0
box -32 -32 32 32
use via_M1_M2_1  NoName_157
timestamp 1647525606
transform 1 0 -256 0 1 0
box -32 -32 32 32
use via_M1_M2_1  NoName_158
timestamp 1647525606
transform 1 0 0 0 1 0
box -32 -32 32 32
use via_M1_M2_1  NoName_159
timestamp 1647525606
transform 1 0 256 0 1 0
box -32 -32 32 32
use via_M1_M2_1  NoName_160
timestamp 1647525606
transform 1 0 512 0 1 0
box -32 -32 32 32
use via_M1_M2_1  NoName_161
timestamp 1647525606
transform 1 0 768 0 1 0
box -32 -32 32 32
use via_M1_M2_1  NoName_162
timestamp 1647525606
transform 1 0 1024 0 1 0
box -32 -32 32 32
use via_M1_M2_1  NoName_163
timestamp 1647525606
transform 1 0 1280 0 1 0
box -32 -32 32 32
use via_M1_M2_1  NoName_164
timestamp 1647525606
transform 1 0 1536 0 1 0
box -32 -32 32 32
use via_M1_M2_1  NoName_165
timestamp 1647525606
transform 1 0 1792 0 1 0
box -32 -32 32 32
use via_M1_M2_1  NoName_166
timestamp 1647525606
transform 1 0 2048 0 1 0
box -32 -32 32 32
use via_M1_M2_1  NoName_167
timestamp 1647525606
transform 1 0 2304 0 1 0
box -32 -32 32 32
use via_M1_M2_1  NoName_168
timestamp 1647525606
transform 1 0 2560 0 1 0
box -32 -32 32 32
use via_M1_M2_1  NoName_169
timestamp 1647525606
transform 1 0 -2432 0 1 -400
box -32 -32 32 32
use via_M1_M2_1  NoName_170
timestamp 1647525606
transform 1 0 -2176 0 1 -400
box -32 -32 32 32
use via_M1_M2_1  NoName_171
timestamp 1647525606
transform 1 0 -1920 0 1 -400
box -32 -32 32 32
use via_M1_M2_1  NoName_172
timestamp 1647525606
transform 1 0 -1664 0 1 -400
box -32 -32 32 32
use via_M1_M2_1  NoName_173
timestamp 1647525606
transform 1 0 -1408 0 1 -400
box -32 -32 32 32
use via_M1_M2_1  NoName_174
timestamp 1647525606
transform 1 0 -1152 0 1 -400
box -32 -32 32 32
use via_M1_M2_1  NoName_175
timestamp 1647525606
transform 1 0 -896 0 1 -400
box -32 -32 32 32
use via_M1_M2_1  NoName_176
timestamp 1647525606
transform 1 0 -640 0 1 -400
box -32 -32 32 32
use via_M1_M2_1  NoName_177
timestamp 1647525606
transform 1 0 -384 0 1 -400
box -32 -32 32 32
use via_M1_M2_1  NoName_178
timestamp 1647525606
transform 1 0 -128 0 1 -400
box -32 -32 32 32
use via_M1_M2_1  NoName_179
timestamp 1647525606
transform 1 0 128 0 1 -400
box -32 -32 32 32
use via_M1_M2_1  NoName_180
timestamp 1647525606
transform 1 0 384 0 1 -400
box -32 -32 32 32
use via_M1_M2_1  NoName_181
timestamp 1647525606
transform 1 0 640 0 1 -400
box -32 -32 32 32
use via_M1_M2_1  NoName_182
timestamp 1647525606
transform 1 0 896 0 1 -400
box -32 -32 32 32
use via_M1_M2_1  NoName_183
timestamp 1647525606
transform 1 0 1152 0 1 -400
box -32 -32 32 32
use via_M1_M2_1  NoName_184
timestamp 1647525606
transform 1 0 1408 0 1 -400
box -32 -32 32 32
use via_M1_M2_1  NoName_185
timestamp 1647525606
transform 1 0 1664 0 1 -400
box -32 -32 32 32
use via_M1_M2_1  NoName_186
timestamp 1647525606
transform 1 0 1920 0 1 -400
box -32 -32 32 32
use via_M1_M2_1  NoName_187
timestamp 1647525606
transform 1 0 2176 0 1 -400
box -32 -32 32 32
use via_M1_M2_1  NoName_188
timestamp 1647525606
transform 1 0 2432 0 1 -400
box -32 -32 32 32
use via_M1_M2_1  NoName_189
timestamp 1647525606
transform 1 0 -2496 0 1 412
box -32 -32 32 32
use via_M1_M2_1  NoName_190
timestamp 1647525606
transform 1 0 -2368 0 1 412
box -32 -32 32 32
use via_M1_M2_1  NoName_191
timestamp 1647525606
transform 1 0 -2240 0 1 412
box -32 -32 32 32
use via_M1_M2_1  NoName_192
timestamp 1647525606
transform 1 0 -2112 0 1 412
box -32 -32 32 32
use via_M1_M2_1  NoName_193
timestamp 1647525606
transform 1 0 -1984 0 1 412
box -32 -32 32 32
use via_M1_M2_1  NoName_194
timestamp 1647525606
transform 1 0 -1854 0 1 412
box -32 -32 32 32
use via_M1_M2_1  NoName_195
timestamp 1647525606
transform 1 0 -1728 0 1 412
box -32 -32 32 32
use via_M1_M2_1  NoName_196
timestamp 1647525606
transform 1 0 -1600 0 1 412
box -32 -32 32 32
use via_M1_M2_1  NoName_197
timestamp 1647525606
transform 1 0 -1472 0 1 412
box -32 -32 32 32
use via_M1_M2_1  NoName_198
timestamp 1647525606
transform 1 0 -1344 0 1 412
box -32 -32 32 32
use via_M1_M2_1  NoName_199
timestamp 1647525606
transform 1 0 -1216 0 1 412
box -32 -32 32 32
use via_M1_M2_1  NoName_200
timestamp 1647525606
transform 1 0 -1088 0 1 412
box -32 -32 32 32
use via_M1_M2_1  NoName_201
timestamp 1647525606
transform 1 0 -960 0 1 412
box -32 -32 32 32
use via_M1_M2_1  NoName_202
timestamp 1647525606
transform 1 0 -832 0 1 412
box -32 -32 32 32
use via_M1_M2_1  NoName_203
timestamp 1647525606
transform 1 0 -704 0 1 412
box -32 -32 32 32
use via_M1_M2_1  NoName_204
timestamp 1647525606
transform 1 0 -576 0 1 412
box -32 -32 32 32
use via_M1_M2_1  NoName_205
timestamp 1647525606
transform 1 0 -448 0 1 412
box -32 -32 32 32
use via_M1_M2_1  NoName_206
timestamp 1647525606
transform 1 0 -320 0 1 412
box -32 -32 32 32
use via_M1_M2_1  NoName_207
timestamp 1647525606
transform 1 0 -192 0 1 412
box -32 -32 32 32
use via_M1_M2_1  NoName_208
timestamp 1647525606
transform 1 0 -64 0 1 412
box -32 -32 32 32
use via_M1_M2_1  NoName_209
timestamp 1647525606
transform 1 0 64 0 1 412
box -32 -32 32 32
use via_M1_M2_1  NoName_210
timestamp 1647525606
transform 1 0 192 0 1 412
box -32 -32 32 32
use via_M1_M2_1  NoName_211
timestamp 1647525606
transform 1 0 320 0 1 412
box -32 -32 32 32
use via_M1_M2_1  NoName_212
timestamp 1647525606
transform 1 0 448 0 1 412
box -32 -32 32 32
use via_M1_M2_1  NoName_213
timestamp 1647525606
transform 1 0 576 0 1 412
box -32 -32 32 32
use via_M1_M2_1  NoName_214
timestamp 1647525606
transform 1 0 704 0 1 412
box -32 -32 32 32
use via_M1_M2_1  NoName_215
timestamp 1647525606
transform 1 0 832 0 1 412
box -32 -32 32 32
use via_M1_M2_1  NoName_216
timestamp 1647525606
transform 1 0 960 0 1 412
box -32 -32 32 32
use via_M1_M2_1  NoName_217
timestamp 1647525606
transform 1 0 1088 0 1 412
box -32 -32 32 32
use via_M1_M2_1  NoName_218
timestamp 1647525606
transform 1 0 1216 0 1 412
box -32 -32 32 32
use via_M1_M2_1  NoName_219
timestamp 1647525606
transform 1 0 1344 0 1 412
box -32 -32 32 32
use via_M1_M2_1  NoName_220
timestamp 1647525606
transform 1 0 1472 0 1 412
box -32 -32 32 32
use via_M1_M2_1  NoName_221
timestamp 1647525606
transform 1 0 1600 0 1 412
box -32 -32 32 32
use via_M1_M2_1  NoName_222
timestamp 1647525606
transform 1 0 1728 0 1 412
box -32 -32 32 32
use via_M1_M2_1  NoName_223
timestamp 1647525606
transform 1 0 1854 0 1 412
box -32 -32 32 32
use via_M1_M2_1  NoName_224
timestamp 1647525606
transform 1 0 1984 0 1 412
box -32 -32 32 32
use via_M1_M2_1  NoName_225
timestamp 1647525606
transform 1 0 2112 0 1 412
box -32 -32 32 32
use via_M1_M2_1  NoName_226
timestamp 1647525606
transform 1 0 2240 0 1 412
box -32 -32 32 32
use via_M1_M2_1  NoName_227
timestamp 1647525606
transform 1 0 2368 0 1 412
box -32 -32 32 32
use via_M1_M2_1  NoName_228
timestamp 1647525606
transform 1 0 2496 0 1 412
box -32 -32 32 32
use XM4_origin  XM4
timestamp 1686232357
transform 1 0 0 0 1 0
box -2727 -534 2727 534
<< end >>
