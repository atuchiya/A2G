magic
tech sky130A
magscale 1 2
timestamp 1686232357
<< checkpaint >>
rect -3987 -1794 3987 1794
<< nwell >>
rect -2727 -534 2727 534
<< pmoslvt >>
rect -2531 -386 -2461 314
rect -2403 -386 -2333 314
rect -2275 -386 -2205 314
rect -2147 -386 -2077 314
rect -2019 -386 -1949 314
rect -1891 -386 -1821 314
rect -1763 -386 -1693 314
rect -1635 -386 -1565 314
rect -1507 -386 -1437 314
rect -1379 -386 -1309 314
rect -1251 -386 -1181 314
rect -1123 -386 -1053 314
rect -995 -386 -925 314
rect -867 -386 -797 314
rect -739 -386 -669 314
rect -611 -386 -541 314
rect -483 -386 -413 314
rect -355 -386 -285 314
rect -227 -386 -157 314
rect -99 -386 -29 314
rect 29 -386 99 314
rect 157 -386 227 314
rect 285 -386 355 314
rect 413 -386 483 314
rect 541 -386 611 314
rect 669 -386 739 314
rect 797 -386 867 314
rect 925 -386 995 314
rect 1053 -386 1123 314
rect 1181 -386 1251 314
rect 1309 -386 1379 314
rect 1437 -386 1507 314
rect 1565 -386 1635 314
rect 1693 -386 1763 314
rect 1821 -386 1891 314
rect 1949 -386 2019 314
rect 2077 -386 2147 314
rect 2205 -386 2275 314
rect 2333 -386 2403 314
rect 2461 -386 2531 314
<< pdiff >>
rect -2589 302 -2531 314
rect -2589 -374 -2577 302
rect -2543 -374 -2531 302
rect -2589 -386 -2531 -374
rect -2461 302 -2403 314
rect -2461 -374 -2449 302
rect -2415 -374 -2403 302
rect -2461 -386 -2403 -374
rect -2333 302 -2275 314
rect -2333 -374 -2321 302
rect -2287 -374 -2275 302
rect -2333 -386 -2275 -374
rect -2205 302 -2147 314
rect -2205 -374 -2193 302
rect -2159 -374 -2147 302
rect -2205 -386 -2147 -374
rect -2077 302 -2019 314
rect -2077 -374 -2065 302
rect -2031 -374 -2019 302
rect -2077 -386 -2019 -374
rect -1949 302 -1891 314
rect -1949 -374 -1937 302
rect -1903 -374 -1891 302
rect -1949 -386 -1891 -374
rect -1821 302 -1763 314
rect -1821 -374 -1809 302
rect -1775 -374 -1763 302
rect -1821 -386 -1763 -374
rect -1693 302 -1635 314
rect -1693 -374 -1681 302
rect -1647 -374 -1635 302
rect -1693 -386 -1635 -374
rect -1565 302 -1507 314
rect -1565 -374 -1553 302
rect -1519 -374 -1507 302
rect -1565 -386 -1507 -374
rect -1437 302 -1379 314
rect -1437 -374 -1425 302
rect -1391 -374 -1379 302
rect -1437 -386 -1379 -374
rect -1309 302 -1251 314
rect -1309 -374 -1297 302
rect -1263 -374 -1251 302
rect -1309 -386 -1251 -374
rect -1181 302 -1123 314
rect -1181 -374 -1169 302
rect -1135 -374 -1123 302
rect -1181 -386 -1123 -374
rect -1053 302 -995 314
rect -1053 -374 -1041 302
rect -1007 -374 -995 302
rect -1053 -386 -995 -374
rect -925 302 -867 314
rect -925 -374 -913 302
rect -879 -374 -867 302
rect -925 -386 -867 -374
rect -797 302 -739 314
rect -797 -374 -785 302
rect -751 -374 -739 302
rect -797 -386 -739 -374
rect -669 302 -611 314
rect -669 -374 -657 302
rect -623 -374 -611 302
rect -669 -386 -611 -374
rect -541 302 -483 314
rect -541 -374 -529 302
rect -495 -374 -483 302
rect -541 -386 -483 -374
rect -413 302 -355 314
rect -413 -374 -401 302
rect -367 -374 -355 302
rect -413 -386 -355 -374
rect -285 302 -227 314
rect -285 -374 -273 302
rect -239 -374 -227 302
rect -285 -386 -227 -374
rect -157 302 -99 314
rect -157 -374 -145 302
rect -111 -374 -99 302
rect -157 -386 -99 -374
rect -29 302 29 314
rect -29 -374 -17 302
rect 17 -374 29 302
rect -29 -386 29 -374
rect 99 302 157 314
rect 99 -374 111 302
rect 145 -374 157 302
rect 99 -386 157 -374
rect 227 302 285 314
rect 227 -374 239 302
rect 273 -374 285 302
rect 227 -386 285 -374
rect 355 302 413 314
rect 355 -374 367 302
rect 401 -374 413 302
rect 355 -386 413 -374
rect 483 302 541 314
rect 483 -374 495 302
rect 529 -374 541 302
rect 483 -386 541 -374
rect 611 302 669 314
rect 611 -374 623 302
rect 657 -374 669 302
rect 611 -386 669 -374
rect 739 302 797 314
rect 739 -374 751 302
rect 785 -374 797 302
rect 739 -386 797 -374
rect 867 302 925 314
rect 867 -374 879 302
rect 913 -374 925 302
rect 867 -386 925 -374
rect 995 302 1053 314
rect 995 -374 1007 302
rect 1041 -374 1053 302
rect 995 -386 1053 -374
rect 1123 302 1181 314
rect 1123 -374 1135 302
rect 1169 -374 1181 302
rect 1123 -386 1181 -374
rect 1251 302 1309 314
rect 1251 -374 1263 302
rect 1297 -374 1309 302
rect 1251 -386 1309 -374
rect 1379 302 1437 314
rect 1379 -374 1391 302
rect 1425 -374 1437 302
rect 1379 -386 1437 -374
rect 1507 302 1565 314
rect 1507 -374 1519 302
rect 1553 -374 1565 302
rect 1507 -386 1565 -374
rect 1635 302 1693 314
rect 1635 -374 1647 302
rect 1681 -374 1693 302
rect 1635 -386 1693 -374
rect 1763 302 1821 314
rect 1763 -374 1775 302
rect 1809 -374 1821 302
rect 1763 -386 1821 -374
rect 1891 302 1949 314
rect 1891 -374 1903 302
rect 1937 -374 1949 302
rect 1891 -386 1949 -374
rect 2019 302 2077 314
rect 2019 -374 2031 302
rect 2065 -374 2077 302
rect 2019 -386 2077 -374
rect 2147 302 2205 314
rect 2147 -374 2159 302
rect 2193 -374 2205 302
rect 2147 -386 2205 -374
rect 2275 302 2333 314
rect 2275 -374 2287 302
rect 2321 -374 2333 302
rect 2275 -386 2333 -374
rect 2403 302 2461 314
rect 2403 -374 2415 302
rect 2449 -374 2461 302
rect 2403 -386 2461 -374
rect 2531 302 2589 314
rect 2531 -374 2543 302
rect 2577 -374 2589 302
rect 2531 -386 2589 -374
<< pdiffc >>
rect -2577 -374 -2543 302
rect -2449 -374 -2415 302
rect -2321 -374 -2287 302
rect -2193 -374 -2159 302
rect -2065 -374 -2031 302
rect -1937 -374 -1903 302
rect -1809 -374 -1775 302
rect -1681 -374 -1647 302
rect -1553 -374 -1519 302
rect -1425 -374 -1391 302
rect -1297 -374 -1263 302
rect -1169 -374 -1135 302
rect -1041 -374 -1007 302
rect -913 -374 -879 302
rect -785 -374 -751 302
rect -657 -374 -623 302
rect -529 -374 -495 302
rect -401 -374 -367 302
rect -273 -374 -239 302
rect -145 -374 -111 302
rect -17 -374 17 302
rect 111 -374 145 302
rect 239 -374 273 302
rect 367 -374 401 302
rect 495 -374 529 302
rect 623 -374 657 302
rect 751 -374 785 302
rect 879 -374 913 302
rect 1007 -374 1041 302
rect 1135 -374 1169 302
rect 1263 -374 1297 302
rect 1391 -374 1425 302
rect 1519 -374 1553 302
rect 1647 -374 1681 302
rect 1775 -374 1809 302
rect 1903 -374 1937 302
rect 2031 -374 2065 302
rect 2159 -374 2193 302
rect 2287 -374 2321 302
rect 2415 -374 2449 302
rect 2543 -374 2577 302
<< nsubdiff >>
rect -2691 464 -2595 498
rect 2595 464 2691 498
rect -2691 401 -2657 464
rect 2657 401 2691 464
rect -2691 -464 -2657 -401
rect 2657 -464 2691 -401
rect -2691 -498 -2595 -464
rect 2595 -498 2691 -464
<< nsubdiffcont >>
rect -2595 464 2595 498
rect -2691 -401 -2657 401
rect 2657 -401 2691 401
rect -2595 -498 2595 -464
<< poly >>
rect -2531 395 -2461 411
rect -2531 361 -2515 395
rect -2477 361 -2461 395
rect -2531 314 -2461 361
rect -2403 395 -2333 411
rect -2403 361 -2387 395
rect -2349 361 -2333 395
rect -2403 314 -2333 361
rect -2275 395 -2205 411
rect -2275 361 -2259 395
rect -2221 361 -2205 395
rect -2275 314 -2205 361
rect -2147 395 -2077 411
rect -2147 361 -2131 395
rect -2093 361 -2077 395
rect -2147 314 -2077 361
rect -2019 395 -1949 411
rect -2019 361 -2003 395
rect -1965 361 -1949 395
rect -2019 314 -1949 361
rect -1891 395 -1821 411
rect -1891 361 -1875 395
rect -1837 361 -1821 395
rect -1891 314 -1821 361
rect -1763 395 -1693 411
rect -1763 361 -1747 395
rect -1709 361 -1693 395
rect -1763 314 -1693 361
rect -1635 395 -1565 411
rect -1635 361 -1619 395
rect -1581 361 -1565 395
rect -1635 314 -1565 361
rect -1507 395 -1437 411
rect -1507 361 -1491 395
rect -1453 361 -1437 395
rect -1507 314 -1437 361
rect -1379 395 -1309 411
rect -1379 361 -1363 395
rect -1325 361 -1309 395
rect -1379 314 -1309 361
rect -1251 395 -1181 411
rect -1251 361 -1235 395
rect -1197 361 -1181 395
rect -1251 314 -1181 361
rect -1123 395 -1053 411
rect -1123 361 -1107 395
rect -1069 361 -1053 395
rect -1123 314 -1053 361
rect -995 395 -925 411
rect -995 361 -979 395
rect -941 361 -925 395
rect -995 314 -925 361
rect -867 395 -797 411
rect -867 361 -851 395
rect -813 361 -797 395
rect -867 314 -797 361
rect -739 395 -669 411
rect -739 361 -723 395
rect -685 361 -669 395
rect -739 314 -669 361
rect -611 395 -541 411
rect -611 361 -595 395
rect -557 361 -541 395
rect -611 314 -541 361
rect -483 395 -413 411
rect -483 361 -467 395
rect -429 361 -413 395
rect -483 314 -413 361
rect -355 395 -285 411
rect -355 361 -339 395
rect -301 361 -285 395
rect -355 314 -285 361
rect -227 395 -157 411
rect -227 361 -211 395
rect -173 361 -157 395
rect -227 314 -157 361
rect -99 395 -29 411
rect -99 361 -83 395
rect -45 361 -29 395
rect -99 314 -29 361
rect 29 395 99 411
rect 29 361 45 395
rect 83 361 99 395
rect 29 314 99 361
rect 157 395 227 411
rect 157 361 173 395
rect 211 361 227 395
rect 157 314 227 361
rect 285 395 355 411
rect 285 361 301 395
rect 339 361 355 395
rect 285 314 355 361
rect 413 395 483 411
rect 413 361 429 395
rect 467 361 483 395
rect 413 314 483 361
rect 541 395 611 411
rect 541 361 557 395
rect 595 361 611 395
rect 541 314 611 361
rect 669 395 739 411
rect 669 361 685 395
rect 723 361 739 395
rect 669 314 739 361
rect 797 395 867 411
rect 797 361 813 395
rect 851 361 867 395
rect 797 314 867 361
rect 925 395 995 411
rect 925 361 941 395
rect 979 361 995 395
rect 925 314 995 361
rect 1053 395 1123 411
rect 1053 361 1069 395
rect 1107 361 1123 395
rect 1053 314 1123 361
rect 1181 395 1251 411
rect 1181 361 1197 395
rect 1235 361 1251 395
rect 1181 314 1251 361
rect 1309 395 1379 411
rect 1309 361 1325 395
rect 1363 361 1379 395
rect 1309 314 1379 361
rect 1437 395 1507 411
rect 1437 361 1453 395
rect 1491 361 1507 395
rect 1437 314 1507 361
rect 1565 395 1635 411
rect 1565 361 1581 395
rect 1619 361 1635 395
rect 1565 314 1635 361
rect 1693 395 1763 411
rect 1693 361 1709 395
rect 1747 361 1763 395
rect 1693 314 1763 361
rect 1821 395 1891 411
rect 1821 361 1837 395
rect 1875 361 1891 395
rect 1821 314 1891 361
rect 1949 395 2019 411
rect 1949 361 1965 395
rect 2003 361 2019 395
rect 1949 314 2019 361
rect 2077 395 2147 411
rect 2077 361 2093 395
rect 2131 361 2147 395
rect 2077 314 2147 361
rect 2205 395 2275 411
rect 2205 361 2221 395
rect 2259 361 2275 395
rect 2205 314 2275 361
rect 2333 395 2403 411
rect 2333 361 2349 395
rect 2387 361 2403 395
rect 2333 314 2403 361
rect 2461 395 2531 411
rect 2461 361 2477 395
rect 2515 361 2531 395
rect 2461 314 2531 361
rect -2531 -412 -2461 -386
rect -2403 -412 -2333 -386
rect -2275 -412 -2205 -386
rect -2147 -412 -2077 -386
rect -2019 -412 -1949 -386
rect -1891 -412 -1821 -386
rect -1763 -412 -1693 -386
rect -1635 -412 -1565 -386
rect -1507 -412 -1437 -386
rect -1379 -412 -1309 -386
rect -1251 -412 -1181 -386
rect -1123 -412 -1053 -386
rect -995 -412 -925 -386
rect -867 -412 -797 -386
rect -739 -412 -669 -386
rect -611 -412 -541 -386
rect -483 -412 -413 -386
rect -355 -412 -285 -386
rect -227 -412 -157 -386
rect -99 -412 -29 -386
rect 29 -412 99 -386
rect 157 -412 227 -386
rect 285 -412 355 -386
rect 413 -412 483 -386
rect 541 -412 611 -386
rect 669 -412 739 -386
rect 797 -412 867 -386
rect 925 -412 995 -386
rect 1053 -412 1123 -386
rect 1181 -412 1251 -386
rect 1309 -412 1379 -386
rect 1437 -412 1507 -386
rect 1565 -412 1635 -386
rect 1693 -412 1763 -386
rect 1821 -412 1891 -386
rect 1949 -412 2019 -386
rect 2077 -412 2147 -386
rect 2205 -412 2275 -386
rect 2333 -412 2403 -386
rect 2461 -412 2531 -386
<< polycont >>
rect -2515 361 -2477 395
rect -2387 361 -2349 395
rect -2259 361 -2221 395
rect -2131 361 -2093 395
rect -2003 361 -1965 395
rect -1875 361 -1837 395
rect -1747 361 -1709 395
rect -1619 361 -1581 395
rect -1491 361 -1453 395
rect -1363 361 -1325 395
rect -1235 361 -1197 395
rect -1107 361 -1069 395
rect -979 361 -941 395
rect -851 361 -813 395
rect -723 361 -685 395
rect -595 361 -557 395
rect -467 361 -429 395
rect -339 361 -301 395
rect -211 361 -173 395
rect -83 361 -45 395
rect 45 361 83 395
rect 173 361 211 395
rect 301 361 339 395
rect 429 361 467 395
rect 557 361 595 395
rect 685 361 723 395
rect 813 361 851 395
rect 941 361 979 395
rect 1069 361 1107 395
rect 1197 361 1235 395
rect 1325 361 1363 395
rect 1453 361 1491 395
rect 1581 361 1619 395
rect 1709 361 1747 395
rect 1837 361 1875 395
rect 1965 361 2003 395
rect 2093 361 2131 395
rect 2221 361 2259 395
rect 2349 361 2387 395
rect 2477 361 2515 395
<< locali >>
rect -2691 464 -2595 498
rect 2595 464 2691 498
rect -2691 401 -2657 464
rect 2657 401 2691 464
rect -2531 361 -2515 395
rect -2477 361 -2461 395
rect -2403 361 -2387 395
rect -2349 361 -2333 395
rect -2275 361 -2259 395
rect -2221 361 -2205 395
rect -2147 361 -2131 395
rect -2093 361 -2077 395
rect -2019 361 -2003 395
rect -1965 361 -1949 395
rect -1891 361 -1875 395
rect -1837 361 -1821 395
rect -1763 361 -1747 395
rect -1709 361 -1693 395
rect -1635 361 -1619 395
rect -1581 361 -1565 395
rect -1507 361 -1491 395
rect -1453 361 -1437 395
rect -1379 361 -1363 395
rect -1325 361 -1309 395
rect -1251 361 -1235 395
rect -1197 361 -1181 395
rect -1123 361 -1107 395
rect -1069 361 -1053 395
rect -995 361 -979 395
rect -941 361 -925 395
rect -867 361 -851 395
rect -813 361 -797 395
rect -739 361 -723 395
rect -685 361 -669 395
rect -611 361 -595 395
rect -557 361 -541 395
rect -483 361 -467 395
rect -429 361 -413 395
rect -355 361 -339 395
rect -301 361 -285 395
rect -227 361 -211 395
rect -173 361 -157 395
rect -99 361 -83 395
rect -45 361 -29 395
rect 29 361 45 395
rect 83 361 99 395
rect 157 361 173 395
rect 211 361 227 395
rect 285 361 301 395
rect 339 361 355 395
rect 413 361 429 395
rect 467 361 483 395
rect 541 361 557 395
rect 595 361 611 395
rect 669 361 685 395
rect 723 361 739 395
rect 797 361 813 395
rect 851 361 867 395
rect 925 361 941 395
rect 979 361 995 395
rect 1053 361 1069 395
rect 1107 361 1123 395
rect 1181 361 1197 395
rect 1235 361 1251 395
rect 1309 361 1325 395
rect 1363 361 1379 395
rect 1437 361 1453 395
rect 1491 361 1507 395
rect 1565 361 1581 395
rect 1619 361 1635 395
rect 1693 361 1709 395
rect 1747 361 1763 395
rect 1821 361 1837 395
rect 1875 361 1891 395
rect 1949 361 1965 395
rect 2003 361 2019 395
rect 2077 361 2093 395
rect 2131 361 2147 395
rect 2205 361 2221 395
rect 2259 361 2275 395
rect 2333 361 2349 395
rect 2387 361 2403 395
rect 2461 361 2477 395
rect 2515 361 2531 395
rect -2577 302 -2543 318
rect -2577 -390 -2543 -374
rect -2449 302 -2415 318
rect -2449 -390 -2415 -374
rect -2321 302 -2287 318
rect -2321 -390 -2287 -374
rect -2193 302 -2159 318
rect -2193 -390 -2159 -374
rect -2065 302 -2031 318
rect -2065 -390 -2031 -374
rect -1937 302 -1903 318
rect -1937 -390 -1903 -374
rect -1809 302 -1775 318
rect -1809 -390 -1775 -374
rect -1681 302 -1647 318
rect -1681 -390 -1647 -374
rect -1553 302 -1519 318
rect -1553 -390 -1519 -374
rect -1425 302 -1391 318
rect -1425 -390 -1391 -374
rect -1297 302 -1263 318
rect -1297 -390 -1263 -374
rect -1169 302 -1135 318
rect -1169 -390 -1135 -374
rect -1041 302 -1007 318
rect -1041 -390 -1007 -374
rect -913 302 -879 318
rect -913 -390 -879 -374
rect -785 302 -751 318
rect -785 -390 -751 -374
rect -657 302 -623 318
rect -657 -390 -623 -374
rect -529 302 -495 318
rect -529 -390 -495 -374
rect -401 302 -367 318
rect -401 -390 -367 -374
rect -273 302 -239 318
rect -273 -390 -239 -374
rect -145 302 -111 318
rect -145 -390 -111 -374
rect -17 302 17 318
rect -17 -390 17 -374
rect 111 302 145 318
rect 111 -390 145 -374
rect 239 302 273 318
rect 239 -390 273 -374
rect 367 302 401 318
rect 367 -390 401 -374
rect 495 302 529 318
rect 495 -390 529 -374
rect 623 302 657 318
rect 623 -390 657 -374
rect 751 302 785 318
rect 751 -390 785 -374
rect 879 302 913 318
rect 879 -390 913 -374
rect 1007 302 1041 318
rect 1007 -390 1041 -374
rect 1135 302 1169 318
rect 1135 -390 1169 -374
rect 1263 302 1297 318
rect 1263 -390 1297 -374
rect 1391 302 1425 318
rect 1391 -390 1425 -374
rect 1519 302 1553 318
rect 1519 -390 1553 -374
rect 1647 302 1681 318
rect 1647 -390 1681 -374
rect 1775 302 1809 318
rect 1775 -390 1809 -374
rect 1903 302 1937 318
rect 1903 -390 1937 -374
rect 2031 302 2065 318
rect 2031 -390 2065 -374
rect 2159 302 2193 318
rect 2159 -390 2193 -374
rect 2287 302 2321 318
rect 2287 -390 2321 -374
rect 2415 302 2449 318
rect 2415 -390 2449 -374
rect 2543 302 2577 318
rect 2543 -390 2577 -374
rect -2691 -464 -2657 -401
rect 2657 -464 2691 -401
rect -2691 -498 -2595 -464
rect 2595 -498 2691 -464
<< viali >>
rect -2515 361 -2477 395
rect -2387 361 -2349 395
rect -2259 361 -2221 395
rect -2131 361 -2093 395
rect -2003 361 -1965 395
rect -1875 361 -1837 395
rect -1747 361 -1709 395
rect -1619 361 -1581 395
rect -1491 361 -1453 395
rect -1363 361 -1325 395
rect -1235 361 -1197 395
rect -1107 361 -1069 395
rect -979 361 -941 395
rect -851 361 -813 395
rect -723 361 -685 395
rect -595 361 -557 395
rect -467 361 -429 395
rect -339 361 -301 395
rect -211 361 -173 395
rect -83 361 -45 395
rect 45 361 83 395
rect 173 361 211 395
rect 301 361 339 395
rect 429 361 467 395
rect 557 361 595 395
rect 685 361 723 395
rect 813 361 851 395
rect 941 361 979 395
rect 1069 361 1107 395
rect 1197 361 1235 395
rect 1325 361 1363 395
rect 1453 361 1491 395
rect 1581 361 1619 395
rect 1709 361 1747 395
rect 1837 361 1875 395
rect 1965 361 2003 395
rect 2093 361 2131 395
rect 2221 361 2259 395
rect 2349 361 2387 395
rect 2477 361 2515 395
rect -2577 -374 -2543 302
rect -2449 -374 -2415 302
rect -2321 -374 -2287 302
rect -2193 -374 -2159 302
rect -2065 -374 -2031 302
rect -1937 -374 -1903 302
rect -1809 -374 -1775 302
rect -1681 -374 -1647 302
rect -1553 -374 -1519 302
rect -1425 -374 -1391 302
rect -1297 -374 -1263 302
rect -1169 -374 -1135 302
rect -1041 -374 -1007 302
rect -913 -374 -879 302
rect -785 -374 -751 302
rect -657 -374 -623 302
rect -529 -374 -495 302
rect -401 -374 -367 302
rect -273 -374 -239 302
rect -145 -374 -111 302
rect -17 -374 17 302
rect 111 -374 145 302
rect 239 -374 273 302
rect 367 -374 401 302
rect 495 -374 529 302
rect 623 -374 657 302
rect 751 -374 785 302
rect 879 -374 913 302
rect 1007 -374 1041 302
rect 1135 -374 1169 302
rect 1263 -374 1297 302
rect 1391 -374 1425 302
rect 1519 -374 1553 302
rect 1647 -374 1681 302
rect 1775 -374 1809 302
rect 1903 -374 1937 302
rect 2031 -374 2065 302
rect 2159 -374 2193 302
rect 2287 -374 2321 302
rect 2415 -374 2449 302
rect 2543 -374 2577 302
<< metal1 >>
rect -2527 395 -2465 401
rect -2527 361 -2515 395
rect -2477 361 -2465 395
rect -2527 355 -2465 361
rect -2399 395 -2337 401
rect -2399 361 -2387 395
rect -2349 361 -2337 395
rect -2399 355 -2337 361
rect -2271 395 -2209 401
rect -2271 361 -2259 395
rect -2221 361 -2209 395
rect -2271 355 -2209 361
rect -2143 395 -2081 401
rect -2143 361 -2131 395
rect -2093 361 -2081 395
rect -2143 355 -2081 361
rect -2015 395 -1953 401
rect -2015 361 -2003 395
rect -1965 361 -1953 395
rect -2015 355 -1953 361
rect -1887 395 -1825 401
rect -1887 361 -1875 395
rect -1837 361 -1825 395
rect -1887 355 -1825 361
rect -1759 395 -1697 401
rect -1759 361 -1747 395
rect -1709 361 -1697 395
rect -1759 355 -1697 361
rect -1631 395 -1569 401
rect -1631 361 -1619 395
rect -1581 361 -1569 395
rect -1631 355 -1569 361
rect -1503 395 -1441 401
rect -1503 361 -1491 395
rect -1453 361 -1441 395
rect -1503 355 -1441 361
rect -1375 395 -1313 401
rect -1375 361 -1363 395
rect -1325 361 -1313 395
rect -1375 355 -1313 361
rect -1247 395 -1185 401
rect -1247 361 -1235 395
rect -1197 361 -1185 395
rect -1247 355 -1185 361
rect -1119 395 -1057 401
rect -1119 361 -1107 395
rect -1069 361 -1057 395
rect -1119 355 -1057 361
rect -991 395 -929 401
rect -991 361 -979 395
rect -941 361 -929 395
rect -991 355 -929 361
rect -863 395 -801 401
rect -863 361 -851 395
rect -813 361 -801 395
rect -863 355 -801 361
rect -735 395 -673 401
rect -735 361 -723 395
rect -685 361 -673 395
rect -735 355 -673 361
rect -607 395 -545 401
rect -607 361 -595 395
rect -557 361 -545 395
rect -607 355 -545 361
rect -479 395 -417 401
rect -479 361 -467 395
rect -429 361 -417 395
rect -479 355 -417 361
rect -351 395 -289 401
rect -351 361 -339 395
rect -301 361 -289 395
rect -351 355 -289 361
rect -223 395 -161 401
rect -223 361 -211 395
rect -173 361 -161 395
rect -223 355 -161 361
rect -95 395 -33 401
rect -95 361 -83 395
rect -45 361 -33 395
rect -95 355 -33 361
rect 33 395 95 401
rect 33 361 45 395
rect 83 361 95 395
rect 33 355 95 361
rect 161 395 223 401
rect 161 361 173 395
rect 211 361 223 395
rect 161 355 223 361
rect 289 395 351 401
rect 289 361 301 395
rect 339 361 351 395
rect 289 355 351 361
rect 417 395 479 401
rect 417 361 429 395
rect 467 361 479 395
rect 417 355 479 361
rect 545 395 607 401
rect 545 361 557 395
rect 595 361 607 395
rect 545 355 607 361
rect 673 395 735 401
rect 673 361 685 395
rect 723 361 735 395
rect 673 355 735 361
rect 801 395 863 401
rect 801 361 813 395
rect 851 361 863 395
rect 801 355 863 361
rect 929 395 991 401
rect 929 361 941 395
rect 979 361 991 395
rect 929 355 991 361
rect 1057 395 1119 401
rect 1057 361 1069 395
rect 1107 361 1119 395
rect 1057 355 1119 361
rect 1185 395 1247 401
rect 1185 361 1197 395
rect 1235 361 1247 395
rect 1185 355 1247 361
rect 1313 395 1375 401
rect 1313 361 1325 395
rect 1363 361 1375 395
rect 1313 355 1375 361
rect 1441 395 1503 401
rect 1441 361 1453 395
rect 1491 361 1503 395
rect 1441 355 1503 361
rect 1569 395 1631 401
rect 1569 361 1581 395
rect 1619 361 1631 395
rect 1569 355 1631 361
rect 1697 395 1759 401
rect 1697 361 1709 395
rect 1747 361 1759 395
rect 1697 355 1759 361
rect 1825 395 1887 401
rect 1825 361 1837 395
rect 1875 361 1887 395
rect 1825 355 1887 361
rect 1953 395 2015 401
rect 1953 361 1965 395
rect 2003 361 2015 395
rect 1953 355 2015 361
rect 2081 395 2143 401
rect 2081 361 2093 395
rect 2131 361 2143 395
rect 2081 355 2143 361
rect 2209 395 2271 401
rect 2209 361 2221 395
rect 2259 361 2271 395
rect 2209 355 2271 361
rect 2337 395 2399 401
rect 2337 361 2349 395
rect 2387 361 2399 395
rect 2337 355 2399 361
rect 2465 395 2527 401
rect 2465 361 2477 395
rect 2515 361 2527 395
rect 2465 355 2527 361
rect -2583 302 -2537 314
rect -2583 -374 -2577 302
rect -2543 -374 -2537 302
rect -2583 -386 -2537 -374
rect -2455 302 -2409 314
rect -2455 -374 -2449 302
rect -2415 -374 -2409 302
rect -2455 -386 -2409 -374
rect -2327 302 -2281 314
rect -2327 -374 -2321 302
rect -2287 -374 -2281 302
rect -2327 -386 -2281 -374
rect -2199 302 -2153 314
rect -2199 -374 -2193 302
rect -2159 -374 -2153 302
rect -2199 -386 -2153 -374
rect -2071 302 -2025 314
rect -2071 -374 -2065 302
rect -2031 -374 -2025 302
rect -2071 -386 -2025 -374
rect -1943 302 -1897 314
rect -1943 -374 -1937 302
rect -1903 -374 -1897 302
rect -1943 -386 -1897 -374
rect -1815 302 -1769 314
rect -1815 -374 -1809 302
rect -1775 -374 -1769 302
rect -1815 -386 -1769 -374
rect -1687 302 -1641 314
rect -1687 -374 -1681 302
rect -1647 -374 -1641 302
rect -1687 -386 -1641 -374
rect -1559 302 -1513 314
rect -1559 -374 -1553 302
rect -1519 -374 -1513 302
rect -1559 -386 -1513 -374
rect -1431 302 -1385 314
rect -1431 -374 -1425 302
rect -1391 -374 -1385 302
rect -1431 -386 -1385 -374
rect -1303 302 -1257 314
rect -1303 -374 -1297 302
rect -1263 -374 -1257 302
rect -1303 -386 -1257 -374
rect -1175 302 -1129 314
rect -1175 -374 -1169 302
rect -1135 -374 -1129 302
rect -1175 -386 -1129 -374
rect -1047 302 -1001 314
rect -1047 -374 -1041 302
rect -1007 -374 -1001 302
rect -1047 -386 -1001 -374
rect -919 302 -873 314
rect -919 -374 -913 302
rect -879 -374 -873 302
rect -919 -386 -873 -374
rect -791 302 -745 314
rect -791 -374 -785 302
rect -751 -374 -745 302
rect -791 -386 -745 -374
rect -663 302 -617 314
rect -663 -374 -657 302
rect -623 -374 -617 302
rect -663 -386 -617 -374
rect -535 302 -489 314
rect -535 -374 -529 302
rect -495 -374 -489 302
rect -535 -386 -489 -374
rect -407 302 -361 314
rect -407 -374 -401 302
rect -367 -374 -361 302
rect -407 -386 -361 -374
rect -279 302 -233 314
rect -279 -374 -273 302
rect -239 -374 -233 302
rect -279 -386 -233 -374
rect -151 302 -105 314
rect -151 -374 -145 302
rect -111 -374 -105 302
rect -151 -386 -105 -374
rect -23 302 23 314
rect -23 -374 -17 302
rect 17 -374 23 302
rect -23 -386 23 -374
rect 105 302 151 314
rect 105 -374 111 302
rect 145 -374 151 302
rect 105 -386 151 -374
rect 233 302 279 314
rect 233 -374 239 302
rect 273 -374 279 302
rect 233 -386 279 -374
rect 361 302 407 314
rect 361 -374 367 302
rect 401 -374 407 302
rect 361 -386 407 -374
rect 489 302 535 314
rect 489 -374 495 302
rect 529 -374 535 302
rect 489 -386 535 -374
rect 617 302 663 314
rect 617 -374 623 302
rect 657 -374 663 302
rect 617 -386 663 -374
rect 745 302 791 314
rect 745 -374 751 302
rect 785 -374 791 302
rect 745 -386 791 -374
rect 873 302 919 314
rect 873 -374 879 302
rect 913 -374 919 302
rect 873 -386 919 -374
rect 1001 302 1047 314
rect 1001 -374 1007 302
rect 1041 -374 1047 302
rect 1001 -386 1047 -374
rect 1129 302 1175 314
rect 1129 -374 1135 302
rect 1169 -374 1175 302
rect 1129 -386 1175 -374
rect 1257 302 1303 314
rect 1257 -374 1263 302
rect 1297 -374 1303 302
rect 1257 -386 1303 -374
rect 1385 302 1431 314
rect 1385 -374 1391 302
rect 1425 -374 1431 302
rect 1385 -386 1431 -374
rect 1513 302 1559 314
rect 1513 -374 1519 302
rect 1553 -374 1559 302
rect 1513 -386 1559 -374
rect 1641 302 1687 314
rect 1641 -374 1647 302
rect 1681 -374 1687 302
rect 1641 -386 1687 -374
rect 1769 302 1815 314
rect 1769 -374 1775 302
rect 1809 -374 1815 302
rect 1769 -386 1815 -374
rect 1897 302 1943 314
rect 1897 -374 1903 302
rect 1937 -374 1943 302
rect 1897 -386 1943 -374
rect 2025 302 2071 314
rect 2025 -374 2031 302
rect 2065 -374 2071 302
rect 2025 -386 2071 -374
rect 2153 302 2199 314
rect 2153 -374 2159 302
rect 2193 -374 2199 302
rect 2153 -386 2199 -374
rect 2281 302 2327 314
rect 2281 -374 2287 302
rect 2321 -374 2327 302
rect 2281 -386 2327 -374
rect 2409 302 2455 314
rect 2409 -374 2415 302
rect 2449 -374 2455 302
rect 2409 -386 2455 -374
rect 2537 302 2583 314
rect 2537 -374 2543 302
rect 2577 -374 2583 302
rect 2537 -386 2583 -374
<< labels >>
flabel metal1 -2496 378 -2496 378 0 FreeSans 240 0 0 0 G
flabel metal1 -2368 378 -2368 378 0 FreeSans 240 0 0 0 G
flabel metal1 -2240 378 -2240 378 0 FreeSans 240 0 0 0 G
flabel metal1 -2112 378 -2112 378 0 FreeSans 240 0 0 0 G
flabel metal1 -1984 378 -1984 378 0 FreeSans 240 0 0 0 G
flabel metal1 -1855 378 -1855 378 0 FreeSans 240 0 0 0 G
flabel metal1 -1728 378 -1728 378 0 FreeSans 240 0 0 0 G
flabel metal1 -1600 378 -1600 378 0 FreeSans 240 0 0 0 G
flabel metal1 -1472 378 -1472 378 0 FreeSans 240 0 0 0 G
flabel metal1 -1344 378 -1344 378 0 FreeSans 240 0 0 0 G
flabel metal1 -1216 378 -1216 378 0 FreeSans 240 0 0 0 G
flabel metal1 -1088 378 -1088 378 0 FreeSans 240 0 0 0 G
flabel metal1 -960 378 -960 378 0 FreeSans 240 0 0 0 G
flabel metal1 -832 378 -832 378 0 FreeSans 240 0 0 0 G
flabel metal1 -704 378 -704 378 0 FreeSans 240 0 0 0 G
flabel metal1 -576 378 -576 378 0 FreeSans 240 0 0 0 G
flabel metal1 -448 378 -448 378 0 FreeSans 240 0 0 0 G
flabel metal1 -320 378 -320 378 0 FreeSans 240 0 0 0 G
flabel metal1 -192 378 -192 378 0 FreeSans 240 0 0 0 G
flabel metal1 -64 378 -64 378 0 FreeSans 240 0 0 0 G
flabel metal1 64 378 64 378 0 FreeSans 240 0 0 0 G
flabel metal1 192 378 192 378 0 FreeSans 240 0 0 0 G
flabel metal1 320 378 320 378 0 FreeSans 240 0 0 0 G
flabel metal1 448 378 448 378 0 FreeSans 240 0 0 0 G
flabel metal1 576 378 576 378 0 FreeSans 240 0 0 0 G
flabel metal1 704 378 704 378 0 FreeSans 240 0 0 0 G
flabel metal1 832 378 832 378 0 FreeSans 240 0 0 0 G
flabel metal1 960 378 960 378 0 FreeSans 240 0 0 0 G
flabel metal1 1088 378 1088 378 0 FreeSans 240 0 0 0 G
flabel metal1 1216 378 1216 378 0 FreeSans 240 0 0 0 G
flabel metal1 1344 378 1344 378 0 FreeSans 240 0 0 0 G
flabel metal1 1472 378 1472 378 0 FreeSans 240 0 0 0 G
flabel metal1 1600 378 1600 378 0 FreeSans 240 0 0 0 G
flabel metal1 1728 378 1728 378 0 FreeSans 240 0 0 0 G
flabel metal1 1855 378 1855 378 0 FreeSans 240 0 0 0 G
flabel metal1 1984 378 1984 378 0 FreeSans 240 0 0 0 G
flabel metal1 2112 378 2112 378 0 FreeSans 240 0 0 0 G
flabel metal1 2240 378 2240 378 0 FreeSans 240 0 0 0 G
flabel metal1 2368 378 2368 378 0 FreeSans 240 0 0 0 G
flabel metal1 2496 378 2496 378 0 FreeSans 240 0 0 0 G
flabel metal1 -2560 -36 -2560 -36 0 FreeSans 240 0 0 0 D
flabel metal1 -2432 -36 -2432 -36 0 FreeSans 240 0 0 0 S
flabel metal1 -2304 -36 -2304 -36 0 FreeSans 240 0 0 0 D
flabel metal1 -2176 -36 -2176 -36 0 FreeSans 240 0 0 0 S
flabel metal1 -2048 -36 -2048 -36 0 FreeSans 240 0 0 0 D
flabel metal1 -1920 -36 -1920 -36 0 FreeSans 240 0 0 0 S
flabel metal1 -1792 -36 -1792 -36 0 FreeSans 240 0 0 0 D
flabel metal1 -1664 -36 -1664 -36 0 FreeSans 240 0 0 0 S
flabel metal1 -1536 -36 -1536 -36 0 FreeSans 240 0 0 0 D
flabel metal1 -1408 -36 -1408 -36 0 FreeSans 240 0 0 0 S
flabel metal1 -1280 -36 -1280 -36 0 FreeSans 240 0 0 0 D
flabel metal1 -1152 -36 -1152 -36 0 FreeSans 240 0 0 0 S
flabel metal1 -1024 -36 -1024 -36 0 FreeSans 240 0 0 0 D
flabel metal1 -896 -36 -896 -36 0 FreeSans 240 0 0 0 S
flabel metal1 -768 -36 -768 -36 0 FreeSans 240 0 0 0 D
flabel metal1 -640 -36 -640 -36 0 FreeSans 240 0 0 0 S
flabel metal1 -512 -36 -512 -36 0 FreeSans 240 0 0 0 D
flabel metal1 -384 -36 -384 -36 0 FreeSans 240 0 0 0 S
flabel metal1 -256 -36 -256 -36 0 FreeSans 240 0 0 0 D
flabel metal1 -128 -36 -128 -36 0 FreeSans 240 0 0 0 S
flabel metal1 0 -36 0 -36 0 FreeSans 240 0 0 0 D
flabel metal1 128 -36 128 -36 0 FreeSans 240 0 0 0 S
flabel metal1 256 -36 256 -36 0 FreeSans 240 0 0 0 D
flabel metal1 384 -36 384 -36 0 FreeSans 240 0 0 0 S
flabel metal1 512 -36 512 -36 0 FreeSans 240 0 0 0 D
flabel metal1 640 -36 640 -36 0 FreeSans 240 0 0 0 S
flabel metal1 768 -36 768 -36 0 FreeSans 240 0 0 0 D
flabel metal1 896 -36 896 -36 0 FreeSans 240 0 0 0 S
flabel metal1 1024 -36 1024 -36 0 FreeSans 240 0 0 0 D
flabel metal1 1152 -36 1152 -36 0 FreeSans 240 0 0 0 S
flabel metal1 1280 -36 1280 -36 0 FreeSans 240 0 0 0 D
flabel metal1 1408 -36 1408 -36 0 FreeSans 240 0 0 0 S
flabel metal1 1536 -36 1536 -36 0 FreeSans 240 0 0 0 D
flabel metal1 1664 -36 1664 -36 0 FreeSans 240 0 0 0 S
flabel metal1 1792 -36 1792 -36 0 FreeSans 240 0 0 0 D
flabel metal1 1920 -36 1920 -36 0 FreeSans 240 0 0 0 S
flabel metal1 2048 -36 2048 -36 0 FreeSans 240 0 0 0 D
flabel metal1 2176 -36 2176 -36 0 FreeSans 240 0 0 0 S
flabel metal1 2304 -36 2304 -36 0 FreeSans 240 0 0 0 D
flabel metal1 2432 -36 2432 -36 0 FreeSans 240 0 0 0 S
flabel metal1 2560 -36 2560 -36 0 FreeSans 240 0 0 0 D
<< properties >>
string FIXED_BBOX -2674 -481 2674 481
<< end >>

