magic
tech sky130A
magscale 1 2
timestamp 1686232357
<< checkpaint >>
rect -3475 -1789 3475 1789
<< pwell >>
rect -2215 -529 2215 529
<< nmoslvt >>
rect -2019 -381 -1949 319
rect -1891 -381 -1821 319
rect -1763 -381 -1693 319
rect -1635 -381 -1565 319
rect -1507 -381 -1437 319
rect -1379 -381 -1309 319
rect -1251 -381 -1181 319
rect -1123 -381 -1053 319
rect -995 -381 -925 319
rect -867 -381 -797 319
rect -739 -381 -669 319
rect -611 -381 -541 319
rect -483 -381 -413 319
rect -355 -381 -285 319
rect -227 -381 -157 319
rect -99 -381 -29 319
rect 29 -381 99 319
rect 157 -381 227 319
rect 285 -381 355 319
rect 413 -381 483 319
rect 541 -381 611 319
rect 669 -381 739 319
rect 797 -381 867 319
rect 925 -381 995 319
rect 1053 -381 1123 319
rect 1181 -381 1251 319
rect 1309 -381 1379 319
rect 1437 -381 1507 319
rect 1565 -381 1635 319
rect 1693 -381 1763 319
rect 1821 -381 1891 319
rect 1949 -381 2019 319
<< ndiff >>
rect -2077 307 -2019 319
rect -2077 -369 -2065 307
rect -2031 -369 -2019 307
rect -2077 -381 -2019 -369
rect -1949 307 -1891 319
rect -1949 -369 -1937 307
rect -1903 -369 -1891 307
rect -1949 -381 -1891 -369
rect -1821 307 -1763 319
rect -1821 -369 -1809 307
rect -1775 -369 -1763 307
rect -1821 -381 -1763 -369
rect -1693 307 -1635 319
rect -1693 -369 -1681 307
rect -1647 -369 -1635 307
rect -1693 -381 -1635 -369
rect -1565 307 -1507 319
rect -1565 -369 -1553 307
rect -1519 -369 -1507 307
rect -1565 -381 -1507 -369
rect -1437 307 -1379 319
rect -1437 -369 -1425 307
rect -1391 -369 -1379 307
rect -1437 -381 -1379 -369
rect -1309 307 -1251 319
rect -1309 -369 -1297 307
rect -1263 -369 -1251 307
rect -1309 -381 -1251 -369
rect -1181 307 -1123 319
rect -1181 -369 -1169 307
rect -1135 -369 -1123 307
rect -1181 -381 -1123 -369
rect -1053 307 -995 319
rect -1053 -369 -1041 307
rect -1007 -369 -995 307
rect -1053 -381 -995 -369
rect -925 307 -867 319
rect -925 -369 -913 307
rect -879 -369 -867 307
rect -925 -381 -867 -369
rect -797 307 -739 319
rect -797 -369 -785 307
rect -751 -369 -739 307
rect -797 -381 -739 -369
rect -669 307 -611 319
rect -669 -369 -657 307
rect -623 -369 -611 307
rect -669 -381 -611 -369
rect -541 307 -483 319
rect -541 -369 -529 307
rect -495 -369 -483 307
rect -541 -381 -483 -369
rect -413 307 -355 319
rect -413 -369 -401 307
rect -367 -369 -355 307
rect -413 -381 -355 -369
rect -285 307 -227 319
rect -285 -369 -273 307
rect -239 -369 -227 307
rect -285 -381 -227 -369
rect -157 307 -99 319
rect -157 -369 -145 307
rect -111 -369 -99 307
rect -157 -381 -99 -369
rect -29 307 29 319
rect -29 -369 -17 307
rect 17 -369 29 307
rect -29 -381 29 -369
rect 99 307 157 319
rect 99 -369 111 307
rect 145 -369 157 307
rect 99 -381 157 -369
rect 227 307 285 319
rect 227 -369 239 307
rect 273 -369 285 307
rect 227 -381 285 -369
rect 355 307 413 319
rect 355 -369 367 307
rect 401 -369 413 307
rect 355 -381 413 -369
rect 483 307 541 319
rect 483 -369 495 307
rect 529 -369 541 307
rect 483 -381 541 -369
rect 611 307 669 319
rect 611 -369 623 307
rect 657 -369 669 307
rect 611 -381 669 -369
rect 739 307 797 319
rect 739 -369 751 307
rect 785 -369 797 307
rect 739 -381 797 -369
rect 867 307 925 319
rect 867 -369 879 307
rect 913 -369 925 307
rect 867 -381 925 -369
rect 995 307 1053 319
rect 995 -369 1007 307
rect 1041 -369 1053 307
rect 995 -381 1053 -369
rect 1123 307 1181 319
rect 1123 -369 1135 307
rect 1169 -369 1181 307
rect 1123 -381 1181 -369
rect 1251 307 1309 319
rect 1251 -369 1263 307
rect 1297 -369 1309 307
rect 1251 -381 1309 -369
rect 1379 307 1437 319
rect 1379 -369 1391 307
rect 1425 -369 1437 307
rect 1379 -381 1437 -369
rect 1507 307 1565 319
rect 1507 -369 1519 307
rect 1553 -369 1565 307
rect 1507 -381 1565 -369
rect 1635 307 1693 319
rect 1635 -369 1647 307
rect 1681 -369 1693 307
rect 1635 -381 1693 -369
rect 1763 307 1821 319
rect 1763 -369 1775 307
rect 1809 -369 1821 307
rect 1763 -381 1821 -369
rect 1891 307 1949 319
rect 1891 -369 1903 307
rect 1937 -369 1949 307
rect 1891 -381 1949 -369
rect 2019 307 2077 319
rect 2019 -369 2031 307
rect 2065 -369 2077 307
rect 2019 -381 2077 -369
<< ndiffc >>
rect -2065 -369 -2031 307
rect -1937 -369 -1903 307
rect -1809 -369 -1775 307
rect -1681 -369 -1647 307
rect -1553 -369 -1519 307
rect -1425 -369 -1391 307
rect -1297 -369 -1263 307
rect -1169 -369 -1135 307
rect -1041 -369 -1007 307
rect -913 -369 -879 307
rect -785 -369 -751 307
rect -657 -369 -623 307
rect -529 -369 -495 307
rect -401 -369 -367 307
rect -273 -369 -239 307
rect -145 -369 -111 307
rect -17 -369 17 307
rect 111 -369 145 307
rect 239 -369 273 307
rect 367 -369 401 307
rect 495 -369 529 307
rect 623 -369 657 307
rect 751 -369 785 307
rect 879 -369 913 307
rect 1007 -369 1041 307
rect 1135 -369 1169 307
rect 1263 -369 1297 307
rect 1391 -369 1425 307
rect 1519 -369 1553 307
rect 1647 -369 1681 307
rect 1775 -369 1809 307
rect 1903 -369 1937 307
rect 2031 -369 2065 307
<< psubdiff >>
rect -2179 459 -2083 493
rect 2083 459 2179 493
rect -2179 397 -2145 459
rect 2145 397 2179 459
rect -2179 -459 -2145 -397
rect 2145 -459 2179 -397
rect -2179 -493 -2083 -459
rect 2083 -493 2179 -459
<< psubdiffcont >>
rect -2083 459 2083 493
rect -2179 -397 -2145 397
rect 2145 -397 2179 397
rect -2083 -493 2083 -459
<< poly >>
rect -2019 391 -1949 407
rect -2019 357 -2003 391
rect -1965 357 -1949 391
rect -2019 319 -1949 357
rect -1891 391 -1821 407
rect -1891 357 -1875 391
rect -1837 357 -1821 391
rect -1891 319 -1821 357
rect -1763 391 -1693 407
rect -1763 357 -1747 391
rect -1709 357 -1693 391
rect -1763 319 -1693 357
rect -1635 391 -1565 407
rect -1635 357 -1619 391
rect -1581 357 -1565 391
rect -1635 319 -1565 357
rect -1507 391 -1437 407
rect -1507 357 -1491 391
rect -1453 357 -1437 391
rect -1507 319 -1437 357
rect -1379 391 -1309 407
rect -1379 357 -1363 391
rect -1325 357 -1309 391
rect -1379 319 -1309 357
rect -1251 391 -1181 407
rect -1251 357 -1235 391
rect -1197 357 -1181 391
rect -1251 319 -1181 357
rect -1123 391 -1053 407
rect -1123 357 -1107 391
rect -1069 357 -1053 391
rect -1123 319 -1053 357
rect -995 391 -925 407
rect -995 357 -979 391
rect -941 357 -925 391
rect -995 319 -925 357
rect -867 391 -797 407
rect -867 357 -851 391
rect -813 357 -797 391
rect -867 319 -797 357
rect -739 391 -669 407
rect -739 357 -723 391
rect -685 357 -669 391
rect -739 319 -669 357
rect -611 391 -541 407
rect -611 357 -595 391
rect -557 357 -541 391
rect -611 319 -541 357
rect -483 391 -413 407
rect -483 357 -467 391
rect -429 357 -413 391
rect -483 319 -413 357
rect -355 391 -285 407
rect -355 357 -339 391
rect -301 357 -285 391
rect -355 319 -285 357
rect -227 391 -157 407
rect -227 357 -211 391
rect -173 357 -157 391
rect -227 319 -157 357
rect -99 391 -29 407
rect -99 357 -83 391
rect -45 357 -29 391
rect -99 319 -29 357
rect 29 391 99 407
rect 29 357 45 391
rect 83 357 99 391
rect 29 319 99 357
rect 157 391 227 407
rect 157 357 173 391
rect 211 357 227 391
rect 157 319 227 357
rect 285 391 355 407
rect 285 357 301 391
rect 339 357 355 391
rect 285 319 355 357
rect 413 391 483 407
rect 413 357 429 391
rect 467 357 483 391
rect 413 319 483 357
rect 541 391 611 407
rect 541 357 557 391
rect 595 357 611 391
rect 541 319 611 357
rect 669 391 739 407
rect 669 357 685 391
rect 723 357 739 391
rect 669 319 739 357
rect 797 391 867 407
rect 797 357 813 391
rect 851 357 867 391
rect 797 319 867 357
rect 925 391 995 407
rect 925 357 941 391
rect 979 357 995 391
rect 925 319 995 357
rect 1053 391 1123 407
rect 1053 357 1069 391
rect 1107 357 1123 391
rect 1053 319 1123 357
rect 1181 391 1251 407
rect 1181 357 1197 391
rect 1235 357 1251 391
rect 1181 319 1251 357
rect 1309 391 1379 407
rect 1309 357 1325 391
rect 1363 357 1379 391
rect 1309 319 1379 357
rect 1437 391 1507 407
rect 1437 357 1453 391
rect 1491 357 1507 391
rect 1437 319 1507 357
rect 1565 391 1635 407
rect 1565 357 1581 391
rect 1619 357 1635 391
rect 1565 319 1635 357
rect 1693 391 1763 407
rect 1693 357 1709 391
rect 1747 357 1763 391
rect 1693 319 1763 357
rect 1821 391 1891 407
rect 1821 357 1837 391
rect 1875 357 1891 391
rect 1821 319 1891 357
rect 1949 391 2019 407
rect 1949 357 1965 391
rect 2003 357 2019 391
rect 1949 319 2019 357
rect -2019 -407 -1949 -381
rect -1891 -407 -1821 -381
rect -1763 -407 -1693 -381
rect -1635 -407 -1565 -381
rect -1507 -407 -1437 -381
rect -1379 -407 -1309 -381
rect -1251 -407 -1181 -381
rect -1123 -407 -1053 -381
rect -995 -407 -925 -381
rect -867 -407 -797 -381
rect -739 -407 -669 -381
rect -611 -407 -541 -381
rect -483 -407 -413 -381
rect -355 -407 -285 -381
rect -227 -407 -157 -381
rect -99 -407 -29 -381
rect 29 -407 99 -381
rect 157 -407 227 -381
rect 285 -407 355 -381
rect 413 -407 483 -381
rect 541 -407 611 -381
rect 669 -407 739 -381
rect 797 -407 867 -381
rect 925 -407 995 -381
rect 1053 -407 1123 -381
rect 1181 -407 1251 -381
rect 1309 -407 1379 -381
rect 1437 -407 1507 -381
rect 1565 -407 1635 -381
rect 1693 -407 1763 -381
rect 1821 -407 1891 -381
rect 1949 -407 2019 -381
<< polycont >>
rect -2003 357 -1965 391
rect -1875 357 -1837 391
rect -1747 357 -1709 391
rect -1619 357 -1581 391
rect -1491 357 -1453 391
rect -1363 357 -1325 391
rect -1235 357 -1197 391
rect -1107 357 -1069 391
rect -979 357 -941 391
rect -851 357 -813 391
rect -723 357 -685 391
rect -595 357 -557 391
rect -467 357 -429 391
rect -339 357 -301 391
rect -211 357 -173 391
rect -83 357 -45 391
rect 45 357 83 391
rect 173 357 211 391
rect 301 357 339 391
rect 429 357 467 391
rect 557 357 595 391
rect 685 357 723 391
rect 813 357 851 391
rect 941 357 979 391
rect 1069 357 1107 391
rect 1197 357 1235 391
rect 1325 357 1363 391
rect 1453 357 1491 391
rect 1581 357 1619 391
rect 1709 357 1747 391
rect 1837 357 1875 391
rect 1965 357 2003 391
<< locali >>
rect -2179 459 -2083 493
rect 2083 459 2179 493
rect -2179 397 -2145 459
rect 2145 397 2179 459
rect -2019 357 -2003 391
rect -1965 357 -1949 391
rect -1891 357 -1875 391
rect -1837 357 -1821 391
rect -1763 357 -1747 391
rect -1709 357 -1693 391
rect -1635 357 -1619 391
rect -1581 357 -1565 391
rect -1507 357 -1491 391
rect -1453 357 -1437 391
rect -1379 357 -1363 391
rect -1325 357 -1309 391
rect -1251 357 -1235 391
rect -1197 357 -1181 391
rect -1123 357 -1107 391
rect -1069 357 -1053 391
rect -995 357 -979 391
rect -941 357 -925 391
rect -867 357 -851 391
rect -813 357 -797 391
rect -739 357 -723 391
rect -685 357 -669 391
rect -611 357 -595 391
rect -557 357 -541 391
rect -483 357 -467 391
rect -429 357 -413 391
rect -355 357 -339 391
rect -301 357 -285 391
rect -227 357 -211 391
rect -173 357 -157 391
rect -99 357 -83 391
rect -45 357 -29 391
rect 29 357 45 391
rect 83 357 99 391
rect 157 357 173 391
rect 211 357 227 391
rect 285 357 301 391
rect 339 357 355 391
rect 413 357 429 391
rect 467 357 483 391
rect 541 357 557 391
rect 595 357 611 391
rect 669 357 685 391
rect 723 357 739 391
rect 797 357 813 391
rect 851 357 867 391
rect 925 357 941 391
rect 979 357 995 391
rect 1053 357 1069 391
rect 1107 357 1123 391
rect 1181 357 1197 391
rect 1235 357 1251 391
rect 1309 357 1325 391
rect 1363 357 1379 391
rect 1437 357 1453 391
rect 1491 357 1507 391
rect 1565 357 1581 391
rect 1619 357 1635 391
rect 1693 357 1709 391
rect 1747 357 1763 391
rect 1821 357 1837 391
rect 1875 357 1891 391
rect 1949 357 1965 391
rect 2003 357 2019 391
rect -2065 307 -2031 323
rect -2065 -385 -2031 -369
rect -1937 307 -1903 323
rect -1937 -385 -1903 -369
rect -1809 307 -1775 323
rect -1809 -385 -1775 -369
rect -1681 307 -1647 323
rect -1681 -385 -1647 -369
rect -1553 307 -1519 323
rect -1553 -385 -1519 -369
rect -1425 307 -1391 323
rect -1425 -385 -1391 -369
rect -1297 307 -1263 323
rect -1297 -385 -1263 -369
rect -1169 307 -1135 323
rect -1169 -385 -1135 -369
rect -1041 307 -1007 323
rect -1041 -385 -1007 -369
rect -913 307 -879 323
rect -913 -385 -879 -369
rect -785 307 -751 323
rect -785 -385 -751 -369
rect -657 307 -623 323
rect -657 -385 -623 -369
rect -529 307 -495 323
rect -529 -385 -495 -369
rect -401 307 -367 323
rect -401 -385 -367 -369
rect -273 307 -239 323
rect -273 -385 -239 -369
rect -145 307 -111 323
rect -145 -385 -111 -369
rect -17 307 17 323
rect -17 -385 17 -369
rect 111 307 145 323
rect 111 -385 145 -369
rect 239 307 273 323
rect 239 -385 273 -369
rect 367 307 401 323
rect 367 -385 401 -369
rect 495 307 529 323
rect 495 -385 529 -369
rect 623 307 657 323
rect 623 -385 657 -369
rect 751 307 785 323
rect 751 -385 785 -369
rect 879 307 913 323
rect 879 -385 913 -369
rect 1007 307 1041 323
rect 1007 -385 1041 -369
rect 1135 307 1169 323
rect 1135 -385 1169 -369
rect 1263 307 1297 323
rect 1263 -385 1297 -369
rect 1391 307 1425 323
rect 1391 -385 1425 -369
rect 1519 307 1553 323
rect 1519 -385 1553 -369
rect 1647 307 1681 323
rect 1647 -385 1681 -369
rect 1775 307 1809 323
rect 1775 -385 1809 -369
rect 1903 307 1937 323
rect 1903 -385 1937 -369
rect 2031 307 2065 323
rect 2031 -385 2065 -369
rect -2179 -459 -2145 -397
rect 2145 -459 2179 -397
rect -2179 -493 -2083 -459
rect 2083 -493 2179 -459
<< viali >>
rect -2003 357 -1965 391
rect -1875 357 -1837 391
rect -1747 357 -1709 391
rect -1619 357 -1581 391
rect -1491 357 -1453 391
rect -1363 357 -1325 391
rect -1235 357 -1197 391
rect -1107 357 -1069 391
rect -979 357 -941 391
rect -851 357 -813 391
rect -723 357 -685 391
rect -595 357 -557 391
rect -467 357 -429 391
rect -339 357 -301 391
rect -211 357 -173 391
rect -83 357 -45 391
rect 45 357 83 391
rect 173 357 211 391
rect 301 357 339 391
rect 429 357 467 391
rect 557 357 595 391
rect 685 357 723 391
rect 813 357 851 391
rect 941 357 979 391
rect 1069 357 1107 391
rect 1197 357 1235 391
rect 1325 357 1363 391
rect 1453 357 1491 391
rect 1581 357 1619 391
rect 1709 357 1747 391
rect 1837 357 1875 391
rect 1965 357 2003 391
rect -2065 -369 -2031 307
rect -1937 -369 -1903 307
rect -1809 -369 -1775 307
rect -1681 -369 -1647 307
rect -1553 -369 -1519 307
rect -1425 -369 -1391 307
rect -1297 -369 -1263 307
rect -1169 -369 -1135 307
rect -1041 -369 -1007 307
rect -913 -369 -879 307
rect -785 -369 -751 307
rect -657 -369 -623 307
rect -529 -369 -495 307
rect -401 -369 -367 307
rect -273 -369 -239 307
rect -145 -369 -111 307
rect -17 -369 17 307
rect 111 -369 145 307
rect 239 -369 273 307
rect 367 -369 401 307
rect 495 -369 529 307
rect 623 -369 657 307
rect 751 -369 785 307
rect 879 -369 913 307
rect 1007 -369 1041 307
rect 1135 -369 1169 307
rect 1263 -369 1297 307
rect 1391 -369 1425 307
rect 1519 -369 1553 307
rect 1647 -369 1681 307
rect 1775 -369 1809 307
rect 1903 -369 1937 307
rect 2031 -369 2065 307
<< metal1 >>
rect -2015 391 -1953 397
rect -2015 357 -2003 391
rect -1965 357 -1953 391
rect -2015 351 -1953 357
rect -1887 391 -1825 397
rect -1887 357 -1875 391
rect -1837 357 -1825 391
rect -1887 351 -1825 357
rect -1759 391 -1697 397
rect -1759 357 -1747 391
rect -1709 357 -1697 391
rect -1759 351 -1697 357
rect -1631 391 -1569 397
rect -1631 357 -1619 391
rect -1581 357 -1569 391
rect -1631 351 -1569 357
rect -1503 391 -1441 397
rect -1503 357 -1491 391
rect -1453 357 -1441 391
rect -1503 351 -1441 357
rect -1375 391 -1313 397
rect -1375 357 -1363 391
rect -1325 357 -1313 391
rect -1375 351 -1313 357
rect -1247 391 -1185 397
rect -1247 357 -1235 391
rect -1197 357 -1185 391
rect -1247 351 -1185 357
rect -1119 391 -1057 397
rect -1119 357 -1107 391
rect -1069 357 -1057 391
rect -1119 351 -1057 357
rect -991 391 -929 397
rect -991 357 -979 391
rect -941 357 -929 391
rect -991 351 -929 357
rect -863 391 -801 397
rect -863 357 -851 391
rect -813 357 -801 391
rect -863 351 -801 357
rect -735 391 -673 397
rect -735 357 -723 391
rect -685 357 -673 391
rect -735 351 -673 357
rect -607 391 -545 397
rect -607 357 -595 391
rect -557 357 -545 391
rect -607 351 -545 357
rect -479 391 -417 397
rect -479 357 -467 391
rect -429 357 -417 391
rect -479 351 -417 357
rect -351 391 -289 397
rect -351 357 -339 391
rect -301 357 -289 391
rect -351 351 -289 357
rect -223 391 -161 397
rect -223 357 -211 391
rect -173 357 -161 391
rect -223 351 -161 357
rect -95 391 -33 397
rect -95 357 -83 391
rect -45 357 -33 391
rect -95 351 -33 357
rect 33 391 95 397
rect 33 357 45 391
rect 83 357 95 391
rect 33 351 95 357
rect 161 391 223 397
rect 161 357 173 391
rect 211 357 223 391
rect 161 351 223 357
rect 289 391 351 397
rect 289 357 301 391
rect 339 357 351 391
rect 289 351 351 357
rect 417 391 479 397
rect 417 357 429 391
rect 467 357 479 391
rect 417 351 479 357
rect 545 391 607 397
rect 545 357 557 391
rect 595 357 607 391
rect 545 351 607 357
rect 673 391 735 397
rect 673 357 685 391
rect 723 357 735 391
rect 673 351 735 357
rect 801 391 863 397
rect 801 357 813 391
rect 851 357 863 391
rect 801 351 863 357
rect 929 391 991 397
rect 929 357 941 391
rect 979 357 991 391
rect 929 351 991 357
rect 1057 391 1119 397
rect 1057 357 1069 391
rect 1107 357 1119 391
rect 1057 351 1119 357
rect 1185 391 1247 397
rect 1185 357 1197 391
rect 1235 357 1247 391
rect 1185 351 1247 357
rect 1313 391 1375 397
rect 1313 357 1325 391
rect 1363 357 1375 391
rect 1313 351 1375 357
rect 1441 391 1503 397
rect 1441 357 1453 391
rect 1491 357 1503 391
rect 1441 351 1503 357
rect 1569 391 1631 397
rect 1569 357 1581 391
rect 1619 357 1631 391
rect 1569 351 1631 357
rect 1697 391 1759 397
rect 1697 357 1709 391
rect 1747 357 1759 391
rect 1697 351 1759 357
rect 1825 391 1887 397
rect 1825 357 1837 391
rect 1875 357 1887 391
rect 1825 351 1887 357
rect 1953 391 2015 397
rect 1953 357 1965 391
rect 2003 357 2015 391
rect 1953 351 2015 357
rect -2071 307 -2025 319
rect -2071 -369 -2065 307
rect -2031 -369 -2025 307
rect -2071 -381 -2025 -369
rect -1943 307 -1897 319
rect -1943 -369 -1937 307
rect -1903 -369 -1897 307
rect -1943 -381 -1897 -369
rect -1815 307 -1769 319
rect -1815 -369 -1809 307
rect -1775 -369 -1769 307
rect -1815 -381 -1769 -369
rect -1687 307 -1641 319
rect -1687 -369 -1681 307
rect -1647 -369 -1641 307
rect -1687 -381 -1641 -369
rect -1559 307 -1513 319
rect -1559 -369 -1553 307
rect -1519 -369 -1513 307
rect -1559 -381 -1513 -369
rect -1431 307 -1385 319
rect -1431 -369 -1425 307
rect -1391 -369 -1385 307
rect -1431 -381 -1385 -369
rect -1303 307 -1257 319
rect -1303 -369 -1297 307
rect -1263 -369 -1257 307
rect -1303 -381 -1257 -369
rect -1175 307 -1129 319
rect -1175 -369 -1169 307
rect -1135 -369 -1129 307
rect -1175 -381 -1129 -369
rect -1047 307 -1001 319
rect -1047 -369 -1041 307
rect -1007 -369 -1001 307
rect -1047 -381 -1001 -369
rect -919 307 -873 319
rect -919 -369 -913 307
rect -879 -369 -873 307
rect -919 -381 -873 -369
rect -791 307 -745 319
rect -791 -369 -785 307
rect -751 -369 -745 307
rect -791 -381 -745 -369
rect -663 307 -617 319
rect -663 -369 -657 307
rect -623 -369 -617 307
rect -663 -381 -617 -369
rect -535 307 -489 319
rect -535 -369 -529 307
rect -495 -369 -489 307
rect -535 -381 -489 -369
rect -407 307 -361 319
rect -407 -369 -401 307
rect -367 -369 -361 307
rect -407 -381 -361 -369
rect -279 307 -233 319
rect -279 -369 -273 307
rect -239 -369 -233 307
rect -279 -381 -233 -369
rect -151 307 -105 319
rect -151 -369 -145 307
rect -111 -369 -105 307
rect -151 -381 -105 -369
rect -23 307 23 319
rect -23 -369 -17 307
rect 17 -369 23 307
rect -23 -381 23 -369
rect 105 307 151 319
rect 105 -369 111 307
rect 145 -369 151 307
rect 105 -381 151 -369
rect 233 307 279 319
rect 233 -369 239 307
rect 273 -369 279 307
rect 233 -381 279 -369
rect 361 307 407 319
rect 361 -369 367 307
rect 401 -369 407 307
rect 361 -381 407 -369
rect 489 307 535 319
rect 489 -369 495 307
rect 529 -369 535 307
rect 489 -381 535 -369
rect 617 307 663 319
rect 617 -369 623 307
rect 657 -369 663 307
rect 617 -381 663 -369
rect 745 307 791 319
rect 745 -369 751 307
rect 785 -369 791 307
rect 745 -381 791 -369
rect 873 307 919 319
rect 873 -369 879 307
rect 913 -369 919 307
rect 873 -381 919 -369
rect 1001 307 1047 319
rect 1001 -369 1007 307
rect 1041 -369 1047 307
rect 1001 -381 1047 -369
rect 1129 307 1175 319
rect 1129 -369 1135 307
rect 1169 -369 1175 307
rect 1129 -381 1175 -369
rect 1257 307 1303 319
rect 1257 -369 1263 307
rect 1297 -369 1303 307
rect 1257 -381 1303 -369
rect 1385 307 1431 319
rect 1385 -369 1391 307
rect 1425 -369 1431 307
rect 1385 -381 1431 -369
rect 1513 307 1559 319
rect 1513 -369 1519 307
rect 1553 -369 1559 307
rect 1513 -381 1559 -369
rect 1641 307 1687 319
rect 1641 -369 1647 307
rect 1681 -369 1687 307
rect 1641 -381 1687 -369
rect 1769 307 1815 319
rect 1769 -369 1775 307
rect 1809 -369 1815 307
rect 1769 -381 1815 -369
rect 1897 307 1943 319
rect 1897 -369 1903 307
rect 1937 -369 1943 307
rect 1897 -381 1943 -369
rect 2025 307 2071 319
rect 2025 -369 2031 307
rect 2065 -369 2071 307
rect 2025 -381 2071 -369
<< labels >>
flabel metal1 -1984 374 -1984 374 0 FreeSans 240 0 0 0 G
flabel metal1 -1855 374 -1855 374 0 FreeSans 240 0 0 0 G
flabel metal1 -1728 374 -1728 374 0 FreeSans 240 0 0 0 G
flabel metal1 -1600 374 -1600 374 0 FreeSans 240 0 0 0 G
flabel metal1 -1472 374 -1472 374 0 FreeSans 240 0 0 0 G
flabel metal1 -1344 374 -1344 374 0 FreeSans 240 0 0 0 G
flabel metal1 -1216 374 -1216 374 0 FreeSans 240 0 0 0 G
flabel metal1 -1088 374 -1088 374 0 FreeSans 240 0 0 0 G
flabel metal1 -960 374 -960 374 0 FreeSans 240 0 0 0 G
flabel metal1 -832 374 -832 374 0 FreeSans 240 0 0 0 G
flabel metal1 -704 374 -704 374 0 FreeSans 240 0 0 0 G
flabel metal1 -576 374 -576 374 0 FreeSans 240 0 0 0 G
flabel metal1 -448 374 -448 374 0 FreeSans 240 0 0 0 G
flabel metal1 -320 374 -320 374 0 FreeSans 240 0 0 0 G
flabel metal1 -192 374 -192 374 0 FreeSans 240 0 0 0 G
flabel metal1 -64 374 -64 374 0 FreeSans 240 0 0 0 G
flabel metal1 64 374 64 374 0 FreeSans 240 0 0 0 G
flabel metal1 192 374 192 374 0 FreeSans 240 0 0 0 G
flabel metal1 320 374 320 374 0 FreeSans 240 0 0 0 G
flabel metal1 448 374 448 374 0 FreeSans 240 0 0 0 G
flabel metal1 576 374 576 374 0 FreeSans 240 0 0 0 G
flabel metal1 704 374 704 374 0 FreeSans 240 0 0 0 G
flabel metal1 832 374 832 374 0 FreeSans 240 0 0 0 G
flabel metal1 960 374 960 374 0 FreeSans 240 0 0 0 G
flabel metal1 1088 374 1088 374 0 FreeSans 240 0 0 0 G
flabel metal1 1216 374 1216 374 0 FreeSans 240 0 0 0 G
flabel metal1 1344 374 1344 374 0 FreeSans 240 0 0 0 G
flabel metal1 1472 374 1472 374 0 FreeSans 240 0 0 0 G
flabel metal1 1600 374 1600 374 0 FreeSans 240 0 0 0 G
flabel metal1 1728 374 1728 374 0 FreeSans 240 0 0 0 G
flabel metal1 1855 374 1855 374 0 FreeSans 240 0 0 0 G
flabel metal1 1984 374 1984 374 0 FreeSans 240 0 0 0 G
flabel metal1 -2048 -31 -2048 -31 0 FreeSans 240 0 0 0 D
flabel metal1 -1920 -31 -1920 -31 0 FreeSans 240 0 0 0 S
flabel metal1 -1792 -31 -1792 -31 0 FreeSans 240 0 0 0 D
flabel metal1 -1664 -31 -1664 -31 0 FreeSans 240 0 0 0 S
flabel metal1 -1536 -31 -1536 -31 0 FreeSans 240 0 0 0 D
flabel metal1 -1408 -31 -1408 -31 0 FreeSans 240 0 0 0 S
flabel metal1 -1280 -31 -1280 -31 0 FreeSans 240 0 0 0 D
flabel metal1 -1152 -31 -1152 -31 0 FreeSans 240 0 0 0 S
flabel metal1 -1024 -31 -1024 -31 0 FreeSans 240 0 0 0 D
flabel metal1 -896 -31 -896 -31 0 FreeSans 240 0 0 0 S
flabel metal1 -768 -31 -768 -31 0 FreeSans 240 0 0 0 D
flabel metal1 -640 -31 -640 -31 0 FreeSans 240 0 0 0 S
flabel metal1 -512 -31 -512 -31 0 FreeSans 240 0 0 0 D
flabel metal1 -384 -31 -384 -31 0 FreeSans 240 0 0 0 S
flabel metal1 -256 -31 -256 -31 0 FreeSans 240 0 0 0 D
flabel metal1 -128 -31 -128 -31 0 FreeSans 240 0 0 0 S
flabel metal1 0 -31 0 -31 0 FreeSans 240 0 0 0 D
flabel metal1 128 -31 128 -31 0 FreeSans 240 0 0 0 S
flabel metal1 256 -31 256 -31 0 FreeSans 240 0 0 0 D
flabel metal1 384 -31 384 -31 0 FreeSans 240 0 0 0 S
flabel metal1 512 -31 512 -31 0 FreeSans 240 0 0 0 D
flabel metal1 640 -31 640 -31 0 FreeSans 240 0 0 0 S
flabel metal1 768 -31 768 -31 0 FreeSans 240 0 0 0 D
flabel metal1 896 -31 896 -31 0 FreeSans 240 0 0 0 S
flabel metal1 1024 -31 1024 -31 0 FreeSans 240 0 0 0 D
flabel metal1 1152 -31 1152 -31 0 FreeSans 240 0 0 0 S
flabel metal1 1280 -31 1280 -31 0 FreeSans 240 0 0 0 D
flabel metal1 1408 -31 1408 -31 0 FreeSans 240 0 0 0 S
flabel metal1 1536 -31 1536 -31 0 FreeSans 240 0 0 0 D
flabel metal1 1664 -31 1664 -31 0 FreeSans 240 0 0 0 S
flabel metal1 1792 -31 1792 -31 0 FreeSans 240 0 0 0 D
flabel metal1 1920 -31 1920 -31 0 FreeSans 240 0 0 0 S
flabel metal1 2048 -31 2048 -31 0 FreeSans 240 0 0 0 D
<< properties >>
string FIXED_BBOX -2162 -476 2162 476
<< end >>

