magic
tech sky130A
magscale 1 2
timestamp 1686266351
<< checkpaint >>
rect -1410 5410 9210 5460
rect -1460 -1410 9260 5410
rect -1410 -1460 9210 -1410
<< viali >>
rect 3060 3534 3094 3568
rect 4704 3534 4738 3568
rect 3060 3462 3094 3496
rect 4704 3462 4738 3496
rect 3060 3390 3094 3424
rect 4704 3390 4738 3424
rect 3060 3318 3094 3352
rect 4704 3318 4738 3352
rect 3060 3246 3094 3280
rect 4704 3246 4738 3280
rect 3060 3174 3094 3208
rect 4704 3174 4738 3208
rect 3060 3102 3094 3136
rect 4704 3102 4738 3136
rect 3060 3030 3094 3064
rect 4704 3030 4738 3064
rect 1860 2514 1894 2548
rect 3504 2514 3538 2548
rect 4260 2514 4294 2548
rect 5904 2514 5938 2548
rect 1860 2442 1894 2476
rect 3504 2442 3538 2476
rect 4260 2442 4294 2476
rect 5904 2442 5938 2476
rect 1860 2370 1894 2404
rect 3504 2370 3538 2404
rect 4260 2370 4294 2404
rect 5904 2370 5938 2404
rect 296 2334 330 2368
rect 1468 2334 1502 2368
rect 6296 2334 6330 2368
rect 7468 2334 7502 2368
rect 1860 2298 1894 2332
rect 3504 2298 3538 2332
rect 4260 2298 4294 2332
rect 5904 2298 5938 2332
rect 296 2262 330 2296
rect 1468 2262 1502 2296
rect 6296 2262 6330 2296
rect 7468 2262 7502 2296
rect 1860 2226 1894 2260
rect 3504 2226 3538 2260
rect 4260 2226 4294 2260
rect 5904 2226 5938 2260
rect 296 2190 330 2224
rect 1468 2190 1502 2224
rect 6296 2190 6330 2224
rect 7468 2190 7502 2224
rect 1860 2154 1894 2188
rect 3504 2154 3538 2188
rect 4260 2154 4294 2188
rect 5904 2154 5938 2188
rect 296 2118 330 2152
rect 1468 2118 1502 2152
rect 6296 2118 6330 2152
rect 7468 2118 7502 2152
rect 1860 2082 1894 2116
rect 3504 2082 3538 2116
rect 4260 2082 4294 2116
rect 5904 2082 5938 2116
rect 296 2046 330 2080
rect 1468 2046 1502 2080
rect 6296 2046 6330 2080
rect 7468 2046 7502 2080
rect 1860 2010 1894 2044
rect 3504 2010 3538 2044
rect 4260 2010 4294 2044
rect 5904 2010 5938 2044
rect 296 1974 330 2008
rect 1468 1974 1502 2008
rect 6296 1974 6330 2008
rect 7468 1974 7502 2008
rect 1860 1938 1894 1972
rect 3504 1938 3538 1972
rect 4260 1938 4294 1972
rect 5904 1938 5938 1972
rect 296 1902 330 1936
rect 1468 1902 1502 1936
rect 6296 1902 6330 1936
rect 7468 1902 7502 1936
rect 1860 1866 1894 1900
rect 3504 1866 3538 1900
rect 4260 1866 4294 1900
rect 5904 1866 5938 1900
rect 296 1830 330 1864
rect 1468 1830 1502 1864
rect 6296 1830 6330 1864
rect 7468 1830 7502 1864
rect 1860 1794 1894 1828
rect 3504 1794 3538 1828
rect 4260 1794 4294 1828
rect 5904 1794 5938 1828
rect 1860 1722 1894 1756
rect 3504 1722 3538 1756
rect 4260 1722 4294 1756
rect 5904 1722 5938 1756
rect 1860 1650 1894 1684
rect 3504 1650 3538 1684
rect 4260 1650 4294 1684
rect 5904 1650 5938 1684
rect 296 1134 330 1168
rect 1468 1134 1502 1168
rect 6296 1134 6330 1168
rect 7468 1134 7502 1168
rect 296 1062 330 1096
rect 1468 1062 1502 1096
rect 6296 1062 6330 1096
rect 7468 1062 7502 1096
rect 296 990 330 1024
rect 1468 990 1502 1024
rect 6296 990 6330 1024
rect 7468 990 7502 1024
rect 296 918 330 952
rect 1468 918 1502 952
rect 1860 934 1894 968
rect 3504 934 3538 968
rect 4260 934 4294 968
rect 5904 934 5938 968
rect 6296 918 6330 952
rect 7468 918 7502 952
rect 296 846 330 880
rect 1468 846 1502 880
rect 1860 862 1894 896
rect 3504 862 3538 896
rect 4260 862 4294 896
rect 5904 862 5938 896
rect 6296 846 6330 880
rect 7468 846 7502 880
rect 296 774 330 808
rect 1468 774 1502 808
rect 1860 790 1894 824
rect 3504 790 3538 824
rect 4260 790 4294 824
rect 5904 790 5938 824
rect 6296 774 6330 808
rect 7468 774 7502 808
rect 296 702 330 736
rect 1468 702 1502 736
rect 1860 718 1894 752
rect 3504 718 3538 752
rect 4260 718 4294 752
rect 5904 718 5938 752
rect 6296 702 6330 736
rect 7468 702 7502 736
rect 296 630 330 664
rect 1468 630 1502 664
rect 1860 646 1894 680
rect 3504 646 3538 680
rect 4260 646 4294 680
rect 5904 646 5938 680
rect 6296 630 6330 664
rect 7468 630 7502 664
rect 1860 574 1894 608
rect 3504 574 3538 608
rect 4260 574 4294 608
rect 5904 574 5938 608
rect 1860 502 1894 536
rect 3504 502 3538 536
rect 4260 502 4294 536
rect 5904 502 5938 536
rect 1860 430 1894 464
rect 3504 430 3538 464
rect 4260 430 4294 464
rect 5904 430 5938 464
<< metal1 >>
rect -150 4150 -50 4200
rect 50 4150 150 4200
rect 250 4150 350 4200
rect 450 4150 550 4200
rect 650 4150 750 4200
rect 850 4150 950 4200
rect 1050 4150 1150 4200
rect 1250 4150 1350 4200
rect 1450 4150 1550 4200
rect 1650 4150 1750 4200
rect 1850 4150 1950 4200
rect 2050 4150 2150 4200
rect 2250 4150 2350 4200
rect 2450 4150 2550 4200
rect 2650 4150 2750 4200
rect 2850 4150 2950 4200
rect 3050 4150 3150 4200
rect 3250 4150 3350 4200
rect 3450 4150 3550 4200
rect 3650 4150 3750 4200
rect 3850 4150 3950 4200
rect 4050 4150 4150 4200
rect 4250 4150 4350 4200
rect 4450 4150 4550 4200
rect 4650 4150 4750 4200
rect 4850 4150 4950 4200
rect 5050 4150 5150 4200
rect 5250 4150 5350 4200
rect 5450 4150 5550 4200
rect 5650 4150 5750 4200
rect 5850 4150 5950 4200
rect 6050 4150 6150 4200
rect 6250 4150 6350 4200
rect 6450 4150 6550 4200
rect 6650 4150 6750 4200
rect 6850 4150 6950 4200
rect 7050 4150 7150 4200
rect 7250 4150 7350 4200
rect 7450 4150 7550 4200
rect 7650 4150 7750 4200
rect 7850 4150 7950 4200
rect -200 4050 8000 4150
rect -150 3950 -50 4050
rect 50 3950 150 4050
rect 250 3950 350 4050
rect 450 3950 550 4050
rect 650 3950 750 4050
rect 850 3950 950 4050
rect 1050 3950 1150 4050
rect 1250 3950 1350 4050
rect 1450 3950 1550 4050
rect 1650 3950 1750 4050
rect 1850 3950 1950 4050
rect 2050 3950 2150 4050
rect 2250 3950 2350 4050
rect 2450 3950 2550 4050
rect 2650 3950 2750 4050
rect 2850 3950 2950 4050
rect 3050 3950 3150 4050
rect 3250 3950 3350 4050
rect 3450 3950 3550 4050
rect 3650 3950 3750 4050
rect 3850 3950 3950 4050
rect 4050 3950 4150 4050
rect 4250 3950 4350 4050
rect 4450 3950 4550 4050
rect 4650 3950 4750 4050
rect 4850 3950 4950 4050
rect 5050 3950 5150 4050
rect 5250 3950 5350 4050
rect 5450 3950 5550 4050
rect 5650 3950 5750 4050
rect 5850 3950 5950 4050
rect 6050 3950 6150 4050
rect 6250 3950 6350 4050
rect 6450 3950 6550 4050
rect 6650 3950 6750 4050
rect 6850 3950 6950 4050
rect 7050 3950 7150 4050
rect 7250 3950 7350 4050
rect 7450 3950 7550 4050
rect 7650 3950 7750 4050
rect 7850 3950 7950 4050
rect -200 3850 8000 3950
rect -150 3750 -50 3850
rect 50 3750 150 3850
rect 250 3750 350 3850
rect 450 3750 550 3850
rect 650 3750 750 3850
rect 850 3750 950 3850
rect 1050 3750 1150 3850
rect 1250 3750 1350 3850
rect 1450 3750 1550 3850
rect 1650 3750 1750 3850
rect 1850 3750 1950 3850
rect 2050 3750 2150 3850
rect 2250 3750 2350 3850
rect 2450 3750 2550 3850
rect 2650 3750 2750 3850
rect 2850 3750 2950 3850
rect 3050 3800 3150 3850
rect 3250 3800 3350 3850
rect 3450 3800 3550 3850
rect 3650 3800 3750 3850
rect 3850 3800 3950 3850
rect 4050 3800 4150 3850
rect 4250 3800 4350 3850
rect 4450 3800 4550 3850
rect 4650 3800 4750 3850
rect 4850 3750 4950 3850
rect 5050 3750 5150 3850
rect 5250 3750 5350 3850
rect 5450 3750 5550 3850
rect 5650 3750 5750 3850
rect 5850 3750 5950 3850
rect 6050 3750 6150 3850
rect 6250 3750 6350 3850
rect 6450 3750 6550 3850
rect 6650 3750 6750 3850
rect 6850 3750 6950 3850
rect 7050 3750 7150 3850
rect 7250 3750 7350 3850
rect 7450 3750 7550 3850
rect 7650 3750 7750 3850
rect 7850 3750 7950 3850
rect -200 3650 3000 3750
rect 4800 3650 8000 3750
rect -150 3550 -50 3650
rect 50 3550 150 3650
rect 250 3550 350 3650
rect 450 3550 550 3650
rect 650 3550 750 3650
rect 850 3550 950 3650
rect 1050 3550 1150 3650
rect 1250 3550 1350 3650
rect 1450 3550 1550 3650
rect 1650 3550 1750 3650
rect 1850 3550 1950 3650
rect 2050 3550 2150 3650
rect 2250 3550 2350 3650
rect 2450 3550 2550 3650
rect 2650 3550 2750 3650
rect 2850 3550 2950 3650
rect 3038 3568 3118 3588
rect -200 3450 3000 3550
rect 3038 3534 3060 3568
rect 3094 3534 3118 3568
rect 3038 3496 3118 3534
rect 3038 3462 3060 3496
rect 3094 3462 3118 3496
rect -150 3350 -50 3450
rect 50 3350 150 3450
rect 250 3350 350 3450
rect 450 3350 550 3450
rect 650 3350 750 3450
rect 850 3350 950 3450
rect 1050 3350 1150 3450
rect 1250 3350 1350 3450
rect 1450 3350 1550 3450
rect 1650 3350 1750 3450
rect 1850 3350 1950 3450
rect 2050 3350 2150 3450
rect 2250 3350 2350 3450
rect 2450 3350 2550 3450
rect 2650 3350 2750 3450
rect 2850 3350 2950 3450
rect 3038 3424 3118 3462
rect 3038 3390 3060 3424
rect 3094 3390 3118 3424
rect 3038 3352 3118 3390
rect -200 3250 3000 3350
rect 3038 3318 3060 3352
rect 3094 3318 3118 3352
rect 3038 3280 3118 3318
rect -150 3150 -50 3250
rect 50 3150 150 3250
rect 250 3150 350 3250
rect 450 3150 550 3250
rect 650 3150 750 3250
rect 850 3150 950 3250
rect 1050 3150 1150 3250
rect 1250 3150 1350 3250
rect 1450 3150 1550 3250
rect 1650 3150 1750 3250
rect 1850 3150 1950 3250
rect 2050 3150 2150 3250
rect 2250 3150 2350 3250
rect 2450 3150 2550 3250
rect 2650 3150 2750 3250
rect 2850 3150 2950 3250
rect 3038 3246 3060 3280
rect 3094 3246 3118 3280
rect 3038 3208 3118 3246
rect 3038 3174 3060 3208
rect 3094 3174 3118 3208
rect -200 3050 3000 3150
rect 3038 3136 3118 3174
rect 3038 3102 3060 3136
rect 3094 3102 3118 3136
rect 3038 3064 3118 3102
rect -150 2950 -50 3050
rect 50 2950 150 3050
rect 250 2950 350 3050
rect 450 2950 550 3050
rect 650 2950 750 3050
rect 850 2950 950 3050
rect 1050 2950 1150 3050
rect 1250 2950 1350 3050
rect 1450 2950 1550 3050
rect 1650 2950 1750 3050
rect 1850 2950 1950 3050
rect 2050 2950 2150 3050
rect 2250 2950 2350 3050
rect 2450 2950 2550 3050
rect 2650 2950 2750 3050
rect 2850 2950 2950 3050
rect 3038 3030 3060 3064
rect 3094 3030 3118 3064
rect 3038 3010 3118 3030
rect 4682 3568 4762 3588
rect 4682 3534 4704 3568
rect 4738 3534 4762 3568
rect 4850 3550 4950 3650
rect 5050 3550 5150 3650
rect 5250 3550 5350 3650
rect 5450 3550 5550 3650
rect 5650 3550 5750 3650
rect 5850 3550 5950 3650
rect 6050 3550 6150 3650
rect 6250 3550 6350 3650
rect 6450 3550 6550 3650
rect 6650 3550 6750 3650
rect 6850 3550 6950 3650
rect 7050 3550 7150 3650
rect 7250 3550 7350 3650
rect 7450 3550 7550 3650
rect 7650 3550 7750 3650
rect 7850 3550 7950 3650
rect 4682 3496 4762 3534
rect 4682 3462 4704 3496
rect 4738 3462 4762 3496
rect 4682 3424 4762 3462
rect 4800 3450 8000 3550
rect 4682 3390 4704 3424
rect 4738 3390 4762 3424
rect 4682 3352 4762 3390
rect 4682 3318 4704 3352
rect 4738 3318 4762 3352
rect 4850 3350 4950 3450
rect 5050 3350 5150 3450
rect 5250 3350 5350 3450
rect 5450 3350 5550 3450
rect 5650 3350 5750 3450
rect 5850 3350 5950 3450
rect 6050 3350 6150 3450
rect 6250 3350 6350 3450
rect 6450 3350 6550 3450
rect 6650 3350 6750 3450
rect 6850 3350 6950 3450
rect 7050 3350 7150 3450
rect 7250 3350 7350 3450
rect 7450 3350 7550 3450
rect 7650 3350 7750 3450
rect 7850 3350 7950 3450
rect 4682 3280 4762 3318
rect 4682 3246 4704 3280
rect 4738 3246 4762 3280
rect 4800 3250 8000 3350
rect 4682 3208 4762 3246
rect 4682 3174 4704 3208
rect 4738 3174 4762 3208
rect 4682 3136 4762 3174
rect 4850 3150 4950 3250
rect 5050 3150 5150 3250
rect 5250 3150 5350 3250
rect 5450 3150 5550 3250
rect 5650 3150 5750 3250
rect 5850 3150 5950 3250
rect 6050 3150 6150 3250
rect 6250 3150 6350 3250
rect 6450 3150 6550 3250
rect 6650 3150 6750 3250
rect 6850 3150 6950 3250
rect 7050 3150 7150 3250
rect 7250 3150 7350 3250
rect 7450 3150 7550 3250
rect 7650 3150 7750 3250
rect 7850 3150 7950 3250
rect 4682 3102 4704 3136
rect 4738 3102 4762 3136
rect 4682 3064 4762 3102
rect 4682 3030 4704 3064
rect 4738 3030 4762 3064
rect 4800 3050 8000 3150
rect 4682 3010 4762 3030
rect 4850 2950 4950 3050
rect 5050 2950 5150 3050
rect 5250 2950 5350 3050
rect 5450 2950 5550 3050
rect 5650 2950 5750 3050
rect 5850 2950 5950 3050
rect 6050 2950 6150 3050
rect 6250 2950 6350 3050
rect 6450 2950 6550 3050
rect 6650 2950 6750 3050
rect 6850 2950 6950 3050
rect 7050 2950 7150 3050
rect 7250 2950 7350 3050
rect 7450 2950 7550 3050
rect 7650 2950 7750 3050
rect 7850 2950 7950 3050
rect -200 2850 3000 2950
rect 4800 2850 8000 2950
rect -150 2750 -50 2850
rect 50 2750 150 2850
rect 250 2750 350 2850
rect 450 2750 550 2850
rect 650 2750 750 2850
rect 850 2750 950 2850
rect 1050 2750 1150 2850
rect 1250 2750 1350 2850
rect 1450 2750 1550 2850
rect 1650 2750 1750 2850
rect 1850 2800 1950 2850
rect 2050 2800 2150 2850
rect 2250 2800 2350 2850
rect 2450 2800 2550 2850
rect 2650 2800 2750 2850
rect 2850 2800 2950 2850
rect 4850 2800 4950 2850
rect 5050 2800 5150 2850
rect 5250 2800 5350 2850
rect 5450 2800 5550 2850
rect 5650 2800 5750 2850
rect 5850 2800 5950 2850
rect 3650 2750 3750 2800
rect 3850 2750 3950 2800
rect 4050 2750 4150 2800
rect 6050 2750 6150 2850
rect 6250 2750 6350 2850
rect 6450 2750 6550 2850
rect 6650 2750 6750 2850
rect 6850 2750 6950 2850
rect 7050 2750 7150 2850
rect 7250 2750 7350 2850
rect 7450 2750 7550 2850
rect 7650 2750 7750 2850
rect 7850 2750 7950 2850
rect -200 2650 1800 2750
rect 3600 2650 4200 2750
rect 6000 2650 8000 2750
rect -150 2550 -50 2650
rect 50 2550 150 2650
rect 250 2600 350 2650
rect 450 2600 550 2650
rect 650 2600 750 2650
rect 850 2600 950 2650
rect 1050 2600 1150 2650
rect 1250 2600 1350 2650
rect 1450 2600 1550 2650
rect 1650 2550 1750 2650
rect -200 2450 200 2550
rect 1600 2450 1800 2550
rect 1838 2548 1918 2568
rect 1838 2514 1860 2548
rect 1894 2514 1918 2548
rect 1838 2476 1918 2514
rect -150 2350 -50 2450
rect 50 2350 150 2450
rect 274 2368 354 2388
rect -200 2250 200 2350
rect 274 2334 296 2368
rect 330 2334 354 2368
rect 274 2296 354 2334
rect 274 2262 296 2296
rect 330 2262 354 2296
rect -150 2150 -50 2250
rect 50 2150 150 2250
rect 274 2224 354 2262
rect 274 2190 296 2224
rect 330 2190 354 2224
rect 274 2152 354 2190
rect -200 2050 200 2150
rect 274 2118 296 2152
rect 330 2118 354 2152
rect 274 2080 354 2118
rect -150 1950 -50 2050
rect 50 1950 150 2050
rect 274 2046 296 2080
rect 330 2046 354 2080
rect 274 2008 354 2046
rect 274 1974 296 2008
rect 330 1974 354 2008
rect -200 1850 200 1950
rect 274 1936 354 1974
rect 274 1902 296 1936
rect 330 1902 354 1936
rect 274 1864 354 1902
rect -150 1750 -50 1850
rect 50 1750 150 1850
rect 274 1830 296 1864
rect 330 1830 354 1864
rect 274 1810 354 1830
rect 1446 2368 1526 2388
rect 1446 2334 1468 2368
rect 1502 2334 1526 2368
rect 1650 2350 1750 2450
rect 1838 2442 1860 2476
rect 1894 2442 1918 2476
rect 1838 2404 1918 2442
rect 1838 2370 1860 2404
rect 1894 2370 1918 2404
rect 1446 2296 1526 2334
rect 1446 2262 1468 2296
rect 1502 2262 1526 2296
rect 1446 2224 1526 2262
rect 1600 2250 1800 2350
rect 1838 2332 1918 2370
rect 1838 2298 1860 2332
rect 1894 2298 1918 2332
rect 1838 2260 1918 2298
rect 1446 2190 1468 2224
rect 1502 2190 1526 2224
rect 1446 2152 1526 2190
rect 1446 2118 1468 2152
rect 1502 2118 1526 2152
rect 1650 2150 1750 2250
rect 1838 2226 1860 2260
rect 1894 2226 1918 2260
rect 1838 2188 1918 2226
rect 1838 2154 1860 2188
rect 1894 2154 1918 2188
rect 1446 2080 1526 2118
rect 1446 2046 1468 2080
rect 1502 2046 1526 2080
rect 1600 2050 1800 2150
rect 1838 2116 1918 2154
rect 1838 2082 1860 2116
rect 1894 2082 1918 2116
rect 1446 2008 1526 2046
rect 1446 1974 1468 2008
rect 1502 1974 1526 2008
rect 1446 1936 1526 1974
rect 1650 1950 1750 2050
rect 1838 2044 1918 2082
rect 1838 2010 1860 2044
rect 1894 2010 1918 2044
rect 1838 1972 1918 2010
rect 1446 1902 1468 1936
rect 1502 1902 1526 1936
rect 1446 1864 1526 1902
rect 1446 1830 1468 1864
rect 1502 1830 1526 1864
rect 1600 1850 1800 1950
rect 1838 1938 1860 1972
rect 1894 1938 1918 1972
rect 1838 1900 1918 1938
rect 1838 1866 1860 1900
rect 1894 1866 1918 1900
rect 1446 1810 1526 1830
rect 1650 1750 1750 1850
rect 1838 1828 1918 1866
rect 1838 1794 1860 1828
rect 1894 1794 1918 1828
rect 1838 1756 1918 1794
rect -200 1650 200 1750
rect 1600 1650 1800 1750
rect 1838 1722 1860 1756
rect 1894 1722 1918 1756
rect 1838 1684 1918 1722
rect 1838 1650 1860 1684
rect 1894 1650 1918 1684
rect -150 1550 -50 1650
rect 50 1550 150 1650
rect 250 1550 350 1600
rect 450 1550 550 1600
rect 650 1550 750 1600
rect 850 1550 950 1600
rect 1050 1550 1150 1600
rect 1250 1550 1350 1600
rect 1450 1550 1550 1600
rect 1650 1550 1750 1650
rect 1838 1630 1918 1650
rect 3482 2548 3560 2568
rect 3650 2550 3750 2650
rect 3850 2550 3950 2650
rect 4050 2550 4150 2650
rect 3482 2514 3504 2548
rect 3538 2514 3560 2548
rect 3482 2476 3560 2514
rect 3482 2442 3504 2476
rect 3538 2442 3560 2476
rect 3600 2450 4200 2550
rect 4238 2548 4318 2568
rect 4238 2514 4260 2548
rect 4294 2514 4318 2548
rect 4238 2476 4318 2514
rect 3482 2404 3560 2442
rect 3482 2370 3504 2404
rect 3538 2370 3560 2404
rect 3482 2332 3560 2370
rect 3650 2350 3750 2450
rect 3850 2350 3950 2450
rect 4050 2350 4150 2450
rect 4238 2442 4260 2476
rect 4294 2442 4318 2476
rect 4238 2404 4318 2442
rect 4238 2370 4260 2404
rect 4294 2370 4318 2404
rect 3482 2298 3504 2332
rect 3538 2298 3560 2332
rect 3482 2260 3560 2298
rect 3482 2226 3504 2260
rect 3538 2226 3560 2260
rect 3600 2250 4200 2350
rect 4238 2332 4318 2370
rect 4238 2298 4260 2332
rect 4294 2298 4318 2332
rect 4238 2260 4318 2298
rect 3482 2188 3560 2226
rect 3482 2154 3504 2188
rect 3538 2154 3560 2188
rect 3482 2116 3560 2154
rect 3650 2150 3750 2250
rect 3850 2150 3950 2250
rect 4050 2150 4150 2250
rect 4238 2226 4260 2260
rect 4294 2226 4318 2260
rect 4238 2188 4318 2226
rect 4238 2154 4260 2188
rect 4294 2154 4318 2188
rect 3482 2082 3504 2116
rect 3538 2082 3560 2116
rect 3482 2044 3560 2082
rect 3600 2050 4200 2150
rect 4238 2116 4318 2154
rect 4238 2082 4260 2116
rect 4294 2082 4318 2116
rect 3482 2010 3504 2044
rect 3538 2010 3560 2044
rect 3482 1972 3560 2010
rect 3482 1938 3504 1972
rect 3538 1938 3560 1972
rect 3650 1950 3750 2050
rect 3850 1950 3950 2050
rect 4050 1950 4150 2050
rect 4238 2044 4318 2082
rect 4238 2010 4260 2044
rect 4294 2010 4318 2044
rect 4238 1972 4318 2010
rect 3482 1900 3560 1938
rect 3482 1866 3504 1900
rect 3538 1866 3560 1900
rect 3482 1828 3560 1866
rect 3600 1850 4200 1950
rect 4238 1938 4260 1972
rect 4294 1938 4318 1972
rect 4238 1900 4318 1938
rect 4238 1866 4260 1900
rect 4294 1866 4318 1900
rect 3482 1794 3504 1828
rect 3538 1794 3560 1828
rect 3482 1756 3560 1794
rect 3482 1722 3504 1756
rect 3538 1722 3560 1756
rect 3650 1750 3750 1850
rect 3850 1750 3950 1850
rect 4050 1750 4150 1850
rect 4238 1828 4318 1866
rect 4238 1794 4260 1828
rect 4294 1794 4318 1828
rect 4238 1756 4318 1794
rect 3482 1684 3560 1722
rect 3482 1650 3504 1684
rect 3538 1650 3560 1684
rect 3600 1650 4200 1750
rect 4238 1722 4260 1756
rect 4294 1722 4318 1756
rect 4238 1684 4318 1722
rect 4238 1650 4260 1684
rect 4294 1650 4318 1684
rect 3482 1630 3560 1650
rect 3650 1550 3750 1650
rect 3850 1550 3950 1650
rect 4050 1550 4150 1650
rect 4238 1630 4318 1650
rect 5882 2548 5962 2568
rect 6050 2550 6150 2650
rect 6250 2600 6350 2650
rect 6450 2600 6550 2650
rect 6650 2600 6750 2650
rect 6850 2600 6950 2650
rect 7050 2600 7150 2650
rect 7250 2600 7350 2650
rect 7450 2600 7550 2650
rect 7650 2550 7750 2650
rect 7850 2550 7950 2650
rect 5882 2514 5904 2548
rect 5938 2514 5962 2548
rect 5882 2476 5962 2514
rect 5882 2442 5904 2476
rect 5938 2442 5962 2476
rect 6000 2450 6200 2550
rect 7600 2450 8000 2550
rect 5882 2404 5962 2442
rect 5882 2370 5904 2404
rect 5938 2370 5962 2404
rect 5882 2332 5962 2370
rect 6050 2350 6150 2450
rect 6274 2368 6354 2388
rect 5882 2298 5904 2332
rect 5938 2298 5962 2332
rect 5882 2260 5962 2298
rect 5882 2226 5904 2260
rect 5938 2226 5962 2260
rect 6000 2250 6200 2350
rect 6274 2334 6296 2368
rect 6330 2334 6354 2368
rect 6274 2296 6354 2334
rect 6274 2262 6296 2296
rect 6330 2262 6354 2296
rect 5882 2188 5962 2226
rect 5882 2154 5904 2188
rect 5938 2154 5962 2188
rect 5882 2116 5962 2154
rect 6050 2150 6150 2250
rect 6274 2224 6354 2262
rect 6274 2190 6296 2224
rect 6330 2190 6354 2224
rect 6274 2152 6354 2190
rect 5882 2082 5904 2116
rect 5938 2082 5962 2116
rect 5882 2044 5962 2082
rect 6000 2050 6200 2150
rect 6274 2118 6296 2152
rect 6330 2118 6354 2152
rect 6274 2080 6354 2118
rect 5882 2010 5904 2044
rect 5938 2010 5962 2044
rect 5882 1972 5962 2010
rect 5882 1938 5904 1972
rect 5938 1938 5962 1972
rect 6050 1950 6150 2050
rect 6274 2046 6296 2080
rect 6330 2046 6354 2080
rect 6274 2008 6354 2046
rect 6274 1974 6296 2008
rect 6330 1974 6354 2008
rect 5882 1900 5962 1938
rect 5882 1866 5904 1900
rect 5938 1866 5962 1900
rect 5882 1828 5962 1866
rect 6000 1850 6200 1950
rect 6274 1936 6354 1974
rect 6274 1902 6296 1936
rect 6330 1902 6354 1936
rect 6274 1864 6354 1902
rect 5882 1794 5904 1828
rect 5938 1794 5962 1828
rect 5882 1756 5962 1794
rect 5882 1722 5904 1756
rect 5938 1722 5962 1756
rect 6050 1750 6150 1850
rect 6274 1830 6296 1864
rect 6330 1830 6354 1864
rect 6274 1810 6354 1830
rect 7444 2368 7526 2388
rect 7444 2334 7468 2368
rect 7502 2334 7526 2368
rect 7650 2350 7750 2450
rect 7850 2350 7950 2450
rect 7444 2296 7526 2334
rect 7444 2262 7468 2296
rect 7502 2262 7526 2296
rect 7444 2224 7526 2262
rect 7600 2250 8000 2350
rect 7444 2190 7468 2224
rect 7502 2190 7526 2224
rect 7444 2152 7526 2190
rect 7444 2118 7468 2152
rect 7502 2118 7526 2152
rect 7650 2150 7750 2250
rect 7850 2150 7950 2250
rect 7444 2080 7526 2118
rect 7444 2046 7468 2080
rect 7502 2046 7526 2080
rect 7600 2050 8000 2150
rect 7444 2008 7526 2046
rect 7444 1974 7468 2008
rect 7502 1974 7526 2008
rect 7444 1936 7526 1974
rect 7650 1950 7750 2050
rect 7850 1950 7950 2050
rect 7444 1902 7468 1936
rect 7502 1902 7526 1936
rect 7444 1864 7526 1902
rect 7444 1830 7468 1864
rect 7502 1830 7526 1864
rect 7600 1850 8000 1950
rect 7444 1810 7526 1830
rect 7650 1750 7750 1850
rect 7850 1750 7950 1850
rect 5882 1684 5962 1722
rect 5882 1650 5904 1684
rect 5938 1650 5962 1684
rect 6000 1650 6200 1750
rect 7600 1650 8000 1750
rect 5882 1630 5962 1650
rect 6050 1550 6150 1650
rect 6250 1550 6350 1600
rect 6450 1550 6550 1600
rect 6650 1550 6750 1600
rect 6850 1550 6950 1600
rect 7050 1550 7150 1600
rect 7250 1550 7350 1600
rect 7450 1550 7550 1600
rect 7650 1550 7750 1650
rect 7850 1550 7950 1650
rect -200 1450 1800 1550
rect -150 1350 -50 1450
rect 50 1350 150 1450
rect 250 1400 350 1450
rect 450 1400 550 1450
rect 650 1400 750 1450
rect 850 1400 950 1450
rect 1050 1400 1150 1450
rect 1250 1400 1350 1450
rect 1450 1400 1550 1450
rect 1650 1350 1750 1450
rect 1850 1350 1950 1400
rect 2050 1350 2150 1550
rect 2250 1350 2350 1550
rect 2450 1350 2550 1550
rect 2650 1350 2750 1550
rect 2850 1350 2950 1550
rect 3050 1350 3150 1550
rect 3250 1350 3350 1550
rect 3600 1450 4200 1550
rect 3450 1350 3550 1400
rect 3650 1350 3750 1450
rect 3850 1350 3950 1450
rect 4050 1350 4150 1450
rect 4250 1350 4350 1400
rect 4450 1350 4550 1550
rect 4650 1350 4750 1550
rect 4850 1350 4950 1550
rect 5050 1350 5150 1550
rect 5250 1350 5350 1550
rect 5450 1350 5550 1550
rect 5650 1350 5750 1550
rect 6000 1450 8000 1550
rect 5850 1350 5950 1400
rect 6050 1350 6150 1450
rect 6250 1400 6350 1450
rect 6450 1400 6550 1450
rect 6650 1400 6750 1450
rect 6850 1400 6950 1450
rect 7050 1400 7150 1450
rect 7250 1400 7350 1450
rect 7450 1400 7550 1450
rect 7650 1350 7750 1450
rect 7850 1350 7950 1450
rect -200 1250 200 1350
rect 1600 1250 6200 1350
rect 7600 1250 8000 1350
rect -150 1150 -50 1250
rect 50 1150 150 1250
rect 274 1168 354 1194
rect 274 1150 296 1168
rect -200 1134 296 1150
rect 330 1134 354 1168
rect -200 1096 354 1134
rect -200 1062 296 1096
rect 330 1062 354 1096
rect -200 1050 354 1062
rect -150 950 -50 1050
rect 50 950 150 1050
rect 274 1024 354 1050
rect 274 990 296 1024
rect 330 990 354 1024
rect 274 952 354 990
rect 274 950 296 952
rect -200 918 296 950
rect 330 918 354 952
rect -200 880 354 918
rect -200 850 296 880
rect -150 750 -50 850
rect 50 750 150 850
rect 274 846 296 850
rect 330 846 354 880
rect 274 808 354 846
rect 274 774 296 808
rect 330 774 354 808
rect 274 750 354 774
rect -200 736 354 750
rect -200 702 296 736
rect 330 702 354 736
rect -200 664 354 702
rect -200 650 296 664
rect -150 550 -50 650
rect 50 550 150 650
rect 274 630 296 650
rect 330 630 354 664
rect 274 606 354 630
rect 1446 1168 1526 1194
rect 1446 1134 1468 1168
rect 1502 1150 1526 1168
rect 1650 1150 1750 1250
rect 1850 1200 1950 1250
rect 1502 1134 1800 1150
rect 1446 1096 1800 1134
rect 1446 1062 1468 1096
rect 1502 1062 1800 1096
rect 1446 1050 1800 1062
rect 2050 1050 2150 1250
rect 2250 1050 2350 1250
rect 2450 1050 2550 1250
rect 2650 1050 2750 1250
rect 2850 1050 2950 1250
rect 3050 1050 3150 1250
rect 3250 1050 3350 1250
rect 3450 1200 3550 1250
rect 3650 1150 3750 1250
rect 3850 1150 3950 1250
rect 4050 1150 4150 1250
rect 4250 1200 4350 1250
rect 3600 1050 4200 1150
rect 4450 1050 4550 1250
rect 4650 1050 4750 1250
rect 4850 1050 4950 1250
rect 5050 1050 5150 1250
rect 5250 1050 5350 1250
rect 5450 1050 5550 1250
rect 5650 1050 5750 1250
rect 5850 1200 5950 1250
rect 6050 1150 6150 1250
rect 6274 1168 6354 1194
rect 6274 1150 6296 1168
rect 6000 1134 6296 1150
rect 6330 1134 6354 1168
rect 6000 1096 6354 1134
rect 6000 1062 6296 1096
rect 6330 1062 6354 1096
rect 6000 1050 6354 1062
rect 1446 1024 1526 1050
rect 1446 990 1468 1024
rect 1502 990 1526 1024
rect 1446 952 1526 990
rect 1446 918 1468 952
rect 1502 950 1526 952
rect 1650 950 1750 1050
rect 1838 968 1918 994
rect 1838 950 1860 968
rect 1502 934 1860 950
rect 1894 934 1918 968
rect 1502 918 1918 934
rect 1446 896 1918 918
rect 1446 880 1860 896
rect 1446 846 1468 880
rect 1502 862 1860 880
rect 1894 862 1918 896
rect 1502 850 1918 862
rect 1502 846 1526 850
rect 1446 808 1526 846
rect 1446 774 1468 808
rect 1502 774 1526 808
rect 1446 750 1526 774
rect 1650 750 1750 850
rect 1838 824 1918 850
rect 1838 790 1860 824
rect 1894 790 1918 824
rect 1838 752 1918 790
rect 1838 750 1860 752
rect 1446 736 1860 750
rect 1446 702 1468 736
rect 1502 718 1860 736
rect 1894 718 1918 752
rect 1502 702 1918 718
rect 1446 680 1918 702
rect 1446 664 1860 680
rect 1446 630 1468 664
rect 1502 650 1860 664
rect 1502 630 1526 650
rect 1446 606 1526 630
rect 1650 550 1750 650
rect 1838 646 1860 650
rect 1894 646 1918 680
rect 1838 608 1918 646
rect 1838 574 1860 608
rect 1894 574 1918 608
rect 1838 550 1918 574
rect -200 450 200 550
rect -150 350 -50 450
rect 50 350 150 450
rect 250 350 350 400
rect 450 350 550 400
rect 650 350 750 400
rect 850 350 950 550
rect 1600 536 1918 550
rect 1600 502 1860 536
rect 1894 502 1918 536
rect 1600 464 1918 502
rect 1600 450 1860 464
rect 1050 350 1150 400
rect 1250 350 1350 400
rect 1450 350 1550 400
rect 1650 350 1750 450
rect 1838 430 1860 450
rect 1894 430 1918 464
rect 1838 404 1918 430
rect 3482 968 3560 994
rect 3482 934 3504 968
rect 3538 950 3560 968
rect 3650 950 3750 1050
rect 3850 950 3950 1050
rect 4050 950 4150 1050
rect 4238 968 4318 994
rect 4238 950 4260 968
rect 3538 934 4260 950
rect 4294 934 4318 968
rect 3482 896 4318 934
rect 3482 862 3504 896
rect 3538 862 4260 896
rect 4294 862 4318 896
rect 3482 850 4318 862
rect 3482 824 3560 850
rect 3482 790 3504 824
rect 3538 790 3560 824
rect 3482 752 3560 790
rect 3482 718 3504 752
rect 3538 750 3560 752
rect 3650 750 3750 850
rect 3850 750 3950 850
rect 4050 750 4150 850
rect 4238 824 4318 850
rect 4238 790 4260 824
rect 4294 790 4318 824
rect 4238 752 4318 790
rect 4238 750 4260 752
rect 3538 718 4260 750
rect 4294 718 4318 752
rect 3482 680 4318 718
rect 3482 646 3504 680
rect 3538 650 4260 680
rect 3538 646 3560 650
rect 3482 608 3560 646
rect 3482 574 3504 608
rect 3538 574 3560 608
rect 3482 550 3560 574
rect 3650 550 3750 650
rect 3850 550 3950 650
rect 4050 550 4150 650
rect 4238 646 4260 650
rect 4294 646 4318 680
rect 4238 608 4318 646
rect 4238 574 4260 608
rect 4294 574 4318 608
rect 4238 550 4318 574
rect 3482 536 4318 550
rect 3482 502 3504 536
rect 3538 502 4260 536
rect 4294 502 4318 536
rect 3482 464 4318 502
rect 3482 430 3504 464
rect 3538 450 4260 464
rect 3538 430 3560 450
rect 3482 404 3560 430
rect 3650 350 3750 450
rect 3850 350 3950 450
rect 4050 350 4150 450
rect 4238 430 4260 450
rect 4294 430 4318 464
rect 4238 404 4318 430
rect 5882 968 5962 994
rect 5882 934 5904 968
rect 5938 950 5962 968
rect 6050 950 6150 1050
rect 6274 1024 6354 1050
rect 6274 990 6296 1024
rect 6330 990 6354 1024
rect 6274 952 6354 990
rect 6274 950 6296 952
rect 5938 934 6296 950
rect 5882 918 6296 934
rect 6330 918 6354 952
rect 5882 896 6354 918
rect 5882 862 5904 896
rect 5938 880 6354 896
rect 5938 862 6296 880
rect 5882 850 6296 862
rect 5882 824 5962 850
rect 5882 790 5904 824
rect 5938 790 5962 824
rect 5882 752 5962 790
rect 5882 718 5904 752
rect 5938 750 5962 752
rect 6050 750 6150 850
rect 6274 846 6296 850
rect 6330 846 6354 880
rect 6274 808 6354 846
rect 6274 774 6296 808
rect 6330 774 6354 808
rect 6274 750 6354 774
rect 5938 736 6354 750
rect 5938 718 6296 736
rect 5882 702 6296 718
rect 6330 702 6354 736
rect 5882 680 6354 702
rect 5882 646 5904 680
rect 5938 664 6354 680
rect 5938 650 6296 664
rect 5938 646 5962 650
rect 5882 608 5962 646
rect 5882 574 5904 608
rect 5938 574 5962 608
rect 5882 550 5962 574
rect 6050 550 6150 650
rect 6274 630 6296 650
rect 6330 630 6354 664
rect 6274 606 6354 630
rect 7444 1168 7526 1194
rect 7444 1134 7468 1168
rect 7502 1150 7526 1168
rect 7650 1150 7750 1250
rect 7850 1150 7950 1250
rect 7502 1134 8000 1150
rect 7444 1096 8000 1134
rect 7444 1062 7468 1096
rect 7502 1062 8000 1096
rect 7444 1050 8000 1062
rect 7444 1024 7526 1050
rect 7444 990 7468 1024
rect 7502 990 7526 1024
rect 7444 952 7526 990
rect 7444 918 7468 952
rect 7502 950 7526 952
rect 7650 950 7750 1050
rect 7850 950 7950 1050
rect 7502 918 8000 950
rect 7444 880 8000 918
rect 7444 846 7468 880
rect 7502 850 8000 880
rect 7502 846 7526 850
rect 7444 808 7526 846
rect 7444 774 7468 808
rect 7502 774 7526 808
rect 7444 750 7526 774
rect 7650 750 7750 850
rect 7850 750 7950 850
rect 7444 736 8000 750
rect 7444 702 7468 736
rect 7502 702 8000 736
rect 7444 664 8000 702
rect 7444 630 7468 664
rect 7502 650 8000 664
rect 7502 630 7526 650
rect 7444 606 7526 630
rect 7650 550 7750 650
rect 7850 550 7950 650
rect 5882 536 6200 550
rect 5882 502 5904 536
rect 5938 502 6200 536
rect 5882 464 6200 502
rect 5882 430 5904 464
rect 5938 450 6200 464
rect 5938 430 5962 450
rect 5882 404 5962 430
rect 6050 350 6150 450
rect 6250 350 6350 400
rect 6450 350 6550 400
rect 6650 350 6750 400
rect 6850 350 6950 550
rect 7600 450 8000 550
rect 7050 350 7150 400
rect 7250 350 7350 400
rect 7450 350 7550 400
rect 7650 350 7750 450
rect 7850 350 7950 450
rect -200 250 1800 350
rect 3600 250 4200 350
rect 6000 250 8000 350
rect -150 150 -50 250
rect 50 150 150 250
rect 250 150 350 250
rect 450 150 550 250
rect 650 150 750 250
rect 850 150 950 250
rect 1050 150 1150 250
rect 1250 150 1350 250
rect 1450 150 1550 250
rect 1650 150 1750 250
rect 1850 150 1950 200
rect 2050 150 2150 200
rect 2250 150 2350 200
rect 2450 150 2550 200
rect 2650 150 2750 200
rect 2850 150 2950 200
rect 3050 150 3150 200
rect 3250 150 3350 200
rect 3450 150 3550 200
rect 3650 150 3750 250
rect 3850 150 3950 250
rect 4050 150 4150 250
rect 4250 150 4350 200
rect 4450 150 4550 200
rect 4650 150 4750 200
rect 4850 150 4950 200
rect 5050 150 5150 200
rect 5250 150 5350 200
rect 5450 150 5550 200
rect 5650 150 5750 200
rect 5850 150 5950 200
rect 6050 150 6150 250
rect 6250 150 6350 250
rect 6450 150 6550 250
rect 6650 150 6750 250
rect 6850 150 6950 250
rect 7050 150 7150 250
rect 7250 150 7350 250
rect 7450 150 7550 250
rect 7650 150 7750 250
rect 7850 150 7950 250
rect -200 50 8000 150
rect -150 -50 -50 50
rect 50 -50 150 50
rect 250 -50 350 50
rect 450 -50 550 50
rect 650 -50 750 50
rect 850 -50 950 50
rect 1050 -50 1150 50
rect 1250 -50 1350 50
rect 1450 -50 1550 50
rect 1650 -50 1750 50
rect 1850 -50 1950 50
rect 2050 -50 2150 50
rect 2250 -50 2350 50
rect 2450 -50 2550 50
rect 2650 -50 2750 50
rect 2850 -50 2950 50
rect 3050 -50 3150 50
rect 3250 -50 3350 50
rect 3450 -50 3550 50
rect 3650 -50 3750 50
rect 3850 -50 3950 50
rect 4050 -50 4150 50
rect 4250 -50 4350 50
rect 4450 -50 4550 50
rect 4650 -50 4750 50
rect 4850 -50 4950 50
rect 5050 -50 5150 50
rect 5250 -50 5350 50
rect 5450 -50 5550 50
rect 5650 -50 5750 50
rect 5850 -50 5950 50
rect 6050 -50 6150 50
rect 6250 -50 6350 50
rect 6450 -50 6550 50
rect 6650 -50 6750 50
rect 6850 -50 6950 50
rect 7050 -50 7150 50
rect 7250 -50 7350 50
rect 7450 -50 7550 50
rect 7650 -50 7750 50
rect 7850 -50 7950 50
rect -200 -150 8000 -50
rect -150 -200 -50 -150
rect 50 -200 150 -150
rect 250 -200 350 -150
rect 450 -200 550 -150
rect 650 -200 750 -150
rect 850 -200 950 -150
rect 1050 -200 1150 -150
rect 1250 -200 1350 -150
rect 1450 -200 1550 -150
rect 1650 -200 1750 -150
rect 1850 -200 1950 -150
rect 2050 -200 2150 -150
rect 2250 -200 2350 -150
rect 2450 -200 2550 -150
rect 2650 -200 2750 -150
rect 2850 -200 2950 -150
rect 3050 -200 3150 -150
rect 3250 -200 3350 -150
rect 3450 -200 3550 -150
rect 3650 -200 3750 -150
rect 3850 -200 3950 -150
rect 4050 -200 4150 -150
rect 4250 -200 4350 -150
rect 4450 -200 4550 -150
rect 4650 -200 4750 -150
rect 4850 -200 4950 -150
rect 5050 -200 5150 -150
rect 5250 -200 5350 -150
rect 5450 -200 5550 -150
rect 5650 -200 5750 -150
rect 5850 -200 5950 -150
rect 6050 -200 6150 -150
rect 6250 -200 6350 -150
rect 6450 -200 6550 -150
rect 6650 -200 6750 -150
rect 6850 -200 6950 -150
rect 7050 -200 7150 -150
rect 7250 -200 7350 -150
rect 7450 -200 7550 -150
rect 7650 -200 7750 -150
rect 7850 -200 7950 -150
<< metal2 >>
rect -150 4150 -50 4200
rect 50 4150 150 4200
rect 250 4150 350 4200
rect 450 4150 550 4200
rect 650 4150 750 4200
rect 850 4150 950 4200
rect 1050 4150 1150 4200
rect 1250 4150 1350 4200
rect 1450 4150 1550 4200
rect 1650 4150 1750 4200
rect 1850 4150 1950 4200
rect 2050 4150 2150 4200
rect 2250 4150 2350 4200
rect 2450 4150 2550 4200
rect 2650 4150 2750 4200
rect 2850 4150 2950 4200
rect 3050 4150 3150 4200
rect 3250 4150 3350 4200
rect 3450 4150 3550 4200
rect 3650 4150 3750 4200
rect 3850 4150 3950 4200
rect 4050 4150 4150 4200
rect 4250 4150 4350 4200
rect 4450 4150 4550 4200
rect 4650 4150 4750 4200
rect 4850 4150 4950 4200
rect 5050 4150 5150 4200
rect 5250 4150 5350 4200
rect 5450 4150 5550 4200
rect 5650 4150 5750 4200
rect 5850 4150 5950 4200
rect 6050 4150 6150 4200
rect 6250 4150 6350 4200
rect 6450 4150 6550 4200
rect 6650 4150 6750 4200
rect 6850 4150 6950 4200
rect 7050 4150 7150 4200
rect 7250 4150 7350 4200
rect 7450 4150 7550 4200
rect 7650 4150 7750 4200
rect 7850 4150 7950 4200
rect -200 4050 8000 4150
rect -150 3950 -50 4050
rect 50 3950 150 4050
rect 250 3950 350 4050
rect 450 3950 550 4050
rect 650 3950 750 4050
rect 850 3950 950 4050
rect 1050 3950 1150 4050
rect 1250 3950 1350 4050
rect 1450 3950 1550 4050
rect 1650 3950 1750 4050
rect 1850 3950 1950 4050
rect 2050 3950 2150 4050
rect 2250 3950 2350 4050
rect 2450 3950 2550 4050
rect 2650 3950 2750 4050
rect 2850 3950 2950 4050
rect 3050 3950 3150 4050
rect 3250 3950 3350 4050
rect 3450 3950 3550 4050
rect 3650 3950 3750 4050
rect 3850 3950 3950 4050
rect 4050 3950 4150 4050
rect 4250 3950 4350 4050
rect 4450 3950 4550 4050
rect 4650 3950 4750 4050
rect 4850 3950 4950 4050
rect 5050 3950 5150 4050
rect 5250 3950 5350 4050
rect 5450 3950 5550 4050
rect 5650 3950 5750 4050
rect 5850 3950 5950 4050
rect 6050 3950 6150 4050
rect 6250 3950 6350 4050
rect 6450 3950 6550 4050
rect 6650 3950 6750 4050
rect 6850 3950 6950 4050
rect 7050 3950 7150 4050
rect 7250 3950 7350 4050
rect 7450 3950 7550 4050
rect 7650 3950 7750 4050
rect 7850 3950 7950 4050
rect -200 3850 8000 3950
rect -150 3750 -50 3850
rect 50 3750 150 3850
rect 250 3750 350 3850
rect 450 3750 550 3850
rect 650 3750 750 3850
rect 850 3750 950 3850
rect 1050 3750 1150 3850
rect 1250 3750 1350 3850
rect 1450 3750 1550 3850
rect 1650 3750 1750 3850
rect 1850 3750 1950 3850
rect 2050 3750 2150 3850
rect 2250 3750 2350 3850
rect 2450 3750 2550 3850
rect 2650 3750 2750 3850
rect 2850 3750 2950 3850
rect 3050 3800 3150 3850
rect -200 3650 3000 3750
rect -150 3550 -50 3650
rect 50 3550 150 3650
rect 250 3550 350 3650
rect 450 3550 550 3650
rect 650 3550 750 3650
rect 850 3550 950 3650
rect 1050 3550 1150 3650
rect 1250 3550 1350 3650
rect 1450 3550 1550 3650
rect 1650 3550 1750 3650
rect 1850 3550 1950 3650
rect 2050 3550 2150 3650
rect 2250 3550 2350 3650
rect 2450 3550 2550 3650
rect 2650 3550 2750 3650
rect 2850 3550 2950 3650
rect 3038 3550 3118 3588
rect -200 3450 3118 3550
rect -150 3350 -50 3450
rect 50 3350 150 3450
rect 250 3350 350 3450
rect 450 3350 550 3450
rect 650 3350 750 3450
rect 850 3350 950 3450
rect 1050 3350 1150 3450
rect 1250 3350 1350 3450
rect 1450 3350 1550 3450
rect 1650 3350 1750 3450
rect 1850 3350 1950 3450
rect 2050 3350 2150 3450
rect 2250 3350 2350 3450
rect 2450 3350 2550 3450
rect 2650 3350 2750 3450
rect 2850 3350 2950 3450
rect 3038 3350 3118 3450
rect 3250 3400 3350 3850
rect 3450 3400 3550 3850
rect 3650 3400 3750 3850
rect 3850 3400 3950 3850
rect 4050 3400 4150 3850
rect 4250 3400 4350 3850
rect 4450 3400 4550 3850
rect 4650 3800 4750 3850
rect 4850 3750 4950 3850
rect 5050 3750 5150 3850
rect 5250 3750 5350 3850
rect 5450 3750 5550 3850
rect 5650 3750 5750 3850
rect 5850 3750 5950 3850
rect 6050 3750 6150 3850
rect 6250 3750 6350 3850
rect 6450 3750 6550 3850
rect 6650 3750 6750 3850
rect 6850 3750 6950 3850
rect 7050 3750 7150 3850
rect 7250 3750 7350 3850
rect 7450 3750 7550 3850
rect 7650 3750 7750 3850
rect 7850 3750 7950 3850
rect 4800 3650 8000 3750
rect 4682 3550 4762 3588
rect 4850 3550 4950 3650
rect 5050 3550 5150 3650
rect 5250 3550 5350 3650
rect 5450 3550 5550 3650
rect 5650 3550 5750 3650
rect 5850 3550 5950 3650
rect 6050 3550 6150 3650
rect 6250 3550 6350 3650
rect 6450 3550 6550 3650
rect 6650 3550 6750 3650
rect 6850 3550 6950 3650
rect 7050 3550 7150 3650
rect 7250 3550 7350 3650
rect 7450 3550 7550 3650
rect 7650 3550 7750 3650
rect 7850 3550 7950 3650
rect 4682 3450 8000 3550
rect -200 3250 3118 3350
rect -150 3150 -50 3250
rect 50 3150 150 3250
rect 250 3150 350 3250
rect 450 3150 550 3250
rect 650 3150 750 3250
rect 850 3150 950 3250
rect 1050 3150 1150 3250
rect 1250 3150 1350 3250
rect 1450 3150 1550 3250
rect 1650 3150 1750 3250
rect 1850 3150 1950 3250
rect 2050 3150 2150 3250
rect 2250 3150 2350 3250
rect 2450 3150 2550 3250
rect 2650 3150 2750 3250
rect 2850 3150 2950 3250
rect 3038 3150 3118 3250
rect -200 3050 3118 3150
rect -150 2950 -50 3050
rect 50 2950 150 3050
rect 250 2950 350 3050
rect 450 2950 550 3050
rect 650 2950 750 3050
rect 850 2950 950 3050
rect 1050 2950 1150 3050
rect 1250 2950 1350 3050
rect 1450 2950 1550 3050
rect 1650 2950 1750 3050
rect 1850 2950 1950 3050
rect 2050 2950 2150 3050
rect 2250 2950 2350 3050
rect 2450 2950 2550 3050
rect 2650 2950 2750 3050
rect 2850 2950 2950 3050
rect 3038 3010 3118 3050
rect 4682 3350 4762 3450
rect 4850 3350 4950 3450
rect 5050 3350 5150 3450
rect 5250 3350 5350 3450
rect 5450 3350 5550 3450
rect 5650 3350 5750 3450
rect 5850 3350 5950 3450
rect 6050 3350 6150 3450
rect 6250 3350 6350 3450
rect 6450 3350 6550 3450
rect 6650 3350 6750 3450
rect 6850 3350 6950 3450
rect 7050 3350 7150 3450
rect 7250 3350 7350 3450
rect 7450 3350 7550 3450
rect 7650 3350 7750 3450
rect 7850 3350 7950 3450
rect 4682 3250 8000 3350
rect 4682 3150 4762 3250
rect 4850 3150 4950 3250
rect 5050 3150 5150 3250
rect 5250 3150 5350 3250
rect 5450 3150 5550 3250
rect 5650 3150 5750 3250
rect 5850 3150 5950 3250
rect 6050 3150 6150 3250
rect 6250 3150 6350 3250
rect 6450 3150 6550 3250
rect 6650 3150 6750 3250
rect 6850 3150 6950 3250
rect 7050 3150 7150 3250
rect 7250 3150 7350 3250
rect 7450 3150 7550 3250
rect 7650 3150 7750 3250
rect 7850 3150 7950 3250
rect 4682 3050 8000 3150
rect 4682 3010 4762 3050
rect 4850 2950 4950 3050
rect 5050 2950 5150 3050
rect 5250 2950 5350 3050
rect 5450 2950 5550 3050
rect 5650 2950 5750 3050
rect 5850 2950 5950 3050
rect 6050 2950 6150 3050
rect 6250 2950 6350 3050
rect 6450 2950 6550 3050
rect 6650 2950 6750 3050
rect 6850 2950 6950 3050
rect 7050 2950 7150 3050
rect 7250 2950 7350 3050
rect 7450 2950 7550 3050
rect 7650 2950 7750 3050
rect 7850 2950 7950 3050
rect -200 2850 3000 2950
rect 4800 2850 8000 2950
rect -150 2750 -50 2850
rect 50 2750 150 2850
rect 250 2750 350 2850
rect 450 2750 550 2850
rect 650 2750 750 2850
rect 850 2750 950 2850
rect 1050 2750 1150 2850
rect 1250 2750 1350 2850
rect 1450 2750 1550 2850
rect 1650 2750 1750 2850
rect 1850 2800 1950 2850
rect 2050 2800 2150 2850
rect 2250 2800 2350 2850
rect 2450 2800 2550 2850
rect 2650 2800 2750 2850
rect 2850 2800 2950 2850
rect 4850 2800 4950 2850
rect 5050 2800 5150 2850
rect 5250 2800 5350 2850
rect 5450 2800 5550 2850
rect 5650 2800 5750 2850
rect 5850 2800 5950 2850
rect 3650 2750 3750 2800
rect 3850 2750 3950 2800
rect 4050 2750 4150 2800
rect 6050 2750 6150 2850
rect 6250 2750 6350 2850
rect 6450 2750 6550 2850
rect 6650 2750 6750 2850
rect 6850 2750 6950 2850
rect 7050 2750 7150 2850
rect 7250 2750 7350 2850
rect 7450 2750 7550 2850
rect 7650 2750 7750 2850
rect 7850 2750 7950 2850
rect -200 2650 1800 2750
rect 3600 2650 4200 2750
rect 6000 2650 8000 2750
rect -150 2550 -50 2650
rect 50 2550 150 2650
rect 250 2600 350 2650
rect 450 2600 550 2650
rect 650 2600 750 2650
rect 850 2600 950 2650
rect 1050 2600 1150 2650
rect 1250 2600 1350 2650
rect 1450 2600 1550 2650
rect 1650 2550 1750 2650
rect 1838 2550 1918 2568
rect -200 2450 200 2550
rect 1600 2450 1918 2550
rect -150 2350 -50 2450
rect 50 2350 150 2450
rect 274 2350 354 2388
rect -200 2250 354 2350
rect -150 2150 -50 2250
rect 50 2150 150 2250
rect 274 2150 354 2250
rect -200 2050 354 2150
rect -150 1950 -50 2050
rect 50 1950 150 2050
rect 274 1950 354 2050
rect -200 1850 354 1950
rect -150 1750 -50 1850
rect 50 1750 150 1850
rect 274 1810 354 1850
rect 1446 2350 1526 2388
rect 1650 2350 1750 2450
rect 1838 2350 1918 2450
rect 1446 2250 1918 2350
rect 1446 2150 1526 2250
rect 1650 2150 1750 2250
rect 1838 2150 1918 2250
rect 1446 2050 1918 2150
rect 1446 1950 1526 2050
rect 1650 1950 1750 2050
rect 1838 1950 1918 2050
rect 1446 1850 1918 1950
rect 1446 1810 1526 1850
rect 1650 1750 1750 1850
rect 1838 1750 1918 1850
rect -200 1650 200 1750
rect 1600 1650 1918 1750
rect -150 1550 -50 1650
rect 50 1550 150 1650
rect 250 1550 350 1600
rect 450 1550 550 1600
rect 650 1550 750 1600
rect 850 1550 950 1600
rect 1050 1550 1150 1600
rect 1250 1550 1350 1600
rect 1450 1550 1550 1600
rect 1650 1550 1750 1650
rect 1838 1630 1918 1650
rect 3482 2550 3560 2568
rect 3650 2550 3750 2650
rect 3850 2550 3950 2650
rect 4050 2550 4150 2650
rect 4238 2550 4318 2568
rect 3482 2450 4318 2550
rect 3482 2350 3560 2450
rect 3650 2350 3750 2450
rect 3850 2350 3950 2450
rect 4050 2350 4150 2450
rect 4238 2350 4318 2450
rect 3482 2250 4318 2350
rect 3482 2150 3560 2250
rect 3650 2150 3750 2250
rect 3850 2150 3950 2250
rect 4050 2150 4150 2250
rect 4238 2150 4318 2250
rect 3482 2050 4318 2150
rect 3482 1950 3560 2050
rect 3650 1950 3750 2050
rect 3850 1950 3950 2050
rect 4050 1950 4150 2050
rect 4238 1950 4318 2050
rect 3482 1850 4318 1950
rect 3482 1750 3560 1850
rect 3650 1750 3750 1850
rect 3850 1750 3950 1850
rect 4050 1750 4150 1850
rect 4238 1750 4318 1850
rect 3482 1650 4318 1750
rect 3482 1630 3560 1650
rect 3650 1550 3750 1650
rect 3850 1550 3950 1650
rect 4050 1550 4150 1650
rect 4238 1630 4318 1650
rect 5882 2550 5962 2568
rect 6050 2550 6150 2650
rect 6250 2600 6350 2650
rect 6450 2600 6550 2650
rect 6650 2600 6750 2650
rect 6850 2600 6950 2650
rect 7050 2600 7150 2650
rect 7250 2600 7350 2650
rect 7450 2600 7550 2650
rect 7650 2550 7750 2650
rect 7850 2550 7950 2650
rect 5882 2450 6200 2550
rect 7600 2450 8000 2550
rect 5882 2350 5962 2450
rect 6050 2350 6150 2450
rect 6274 2350 6354 2388
rect 5882 2250 6354 2350
rect 5882 2150 5962 2250
rect 6050 2150 6150 2250
rect 6274 2150 6354 2250
rect 5882 2050 6354 2150
rect 5882 1950 5962 2050
rect 6050 1950 6150 2050
rect 6274 1950 6354 2050
rect 5882 1850 6354 1950
rect 5882 1750 5962 1850
rect 6050 1750 6150 1850
rect 6274 1810 6354 1850
rect 7444 2350 7526 2388
rect 7650 2350 7750 2450
rect 7850 2350 7950 2450
rect 7444 2250 8000 2350
rect 7444 2150 7526 2250
rect 7650 2150 7750 2250
rect 7850 2150 7950 2250
rect 7444 2050 8000 2150
rect 7444 1950 7526 2050
rect 7650 1950 7750 2050
rect 7850 1950 7950 2050
rect 7444 1850 8000 1950
rect 7444 1810 7526 1850
rect 7650 1750 7750 1850
rect 7850 1750 7950 1850
rect 5882 1650 6200 1750
rect 7600 1650 8000 1750
rect 5882 1630 5962 1650
rect 6050 1550 6150 1650
rect 6250 1550 6350 1600
rect 6450 1550 6550 1600
rect 6650 1550 6750 1600
rect 6850 1550 6950 1600
rect 7050 1550 7150 1600
rect 7250 1550 7350 1600
rect 7450 1550 7550 1600
rect 7650 1550 7750 1650
rect 7850 1550 7950 1650
rect -200 1450 1800 1550
rect 3600 1450 4200 1550
rect 6000 1450 8000 1550
rect -150 1350 -50 1450
rect 50 1350 150 1450
rect 250 1400 350 1450
rect 450 1400 550 1450
rect 650 1400 750 1450
rect 850 1400 950 1450
rect 1050 1400 1150 1450
rect 1250 1400 1350 1450
rect 1450 1400 1550 1450
rect 1650 1350 1750 1450
rect 1850 1350 1950 1400
rect 2050 1350 2150 1400
rect 2250 1350 2350 1400
rect 2450 1350 2550 1400
rect 2650 1350 2750 1400
rect 2850 1350 2950 1400
rect 3050 1350 3150 1400
rect 3250 1350 3350 1400
rect 3450 1350 3550 1400
rect 3650 1350 3750 1450
rect 3850 1350 3950 1450
rect 4050 1350 4150 1450
rect 4250 1350 4350 1400
rect 4450 1350 4550 1400
rect 4650 1350 4750 1400
rect 4850 1350 4950 1400
rect 5050 1350 5150 1400
rect 5250 1350 5350 1400
rect 5450 1350 5550 1400
rect 5650 1350 5750 1400
rect 5850 1350 5950 1400
rect 6050 1350 6150 1450
rect 6250 1400 6350 1450
rect 6450 1400 6550 1450
rect 6650 1400 6750 1450
rect 6850 1400 6950 1450
rect 7050 1400 7150 1450
rect 7250 1400 7350 1450
rect 7450 1400 7550 1450
rect 7650 1350 7750 1450
rect 7850 1350 7950 1450
rect -200 1250 200 1350
rect 1600 1250 6200 1350
rect 7600 1250 8000 1350
rect -150 1150 -50 1250
rect 50 1150 150 1250
rect 1650 1150 1750 1250
rect 1850 1200 1950 1250
rect -200 1050 200 1150
rect 1600 1050 1800 1150
rect -150 950 -50 1050
rect 50 950 150 1050
rect 1650 950 1750 1050
rect -200 850 200 950
rect 1600 850 1800 950
rect -150 750 -50 850
rect 50 750 150 850
rect 1650 750 1750 850
rect 2050 800 2150 1250
rect 2250 800 2350 1250
rect 2450 800 2550 1250
rect 2650 800 2750 1250
rect 2850 800 2950 1250
rect 3050 800 3150 1250
rect 3250 800 3350 1250
rect 3450 1200 3550 1250
rect 3650 1150 3750 1250
rect 3850 1150 3950 1250
rect 4050 1150 4150 1250
rect 4250 1200 4350 1250
rect 3600 1050 4200 1150
rect 3650 950 3750 1050
rect 3850 950 3950 1050
rect 4050 950 4150 1050
rect 3600 850 4200 950
rect 3650 750 3750 850
rect 3850 750 3950 850
rect 4050 750 4150 850
rect 4450 800 4550 1250
rect 4650 800 4750 1250
rect 4850 800 4950 1250
rect 5050 800 5150 1250
rect 5250 800 5350 1250
rect 5450 800 5550 1250
rect 5650 800 5750 1250
rect 5850 1200 5950 1250
rect 6050 1150 6150 1250
rect 7650 1150 7750 1250
rect 7850 1150 7950 1250
rect 6000 1050 6200 1150
rect 7600 1050 8000 1150
rect 6050 950 6150 1050
rect 7650 950 7750 1050
rect 7850 950 7950 1050
rect 6000 850 6200 950
rect 7600 850 8000 950
rect 6050 750 6150 850
rect 7650 750 7750 850
rect 7850 750 7950 850
rect -200 650 200 750
rect -150 550 -50 650
rect 50 550 150 650
rect -200 450 200 550
rect 850 500 950 700
rect 1600 650 1800 750
rect 3600 650 4200 750
rect 6000 650 6200 750
rect 1650 550 1750 650
rect 3650 550 3750 650
rect 3850 550 3950 650
rect 4050 550 4150 650
rect 6050 550 6150 650
rect 1600 450 1800 550
rect 3600 450 4200 550
rect 6000 450 6200 550
rect 6850 500 6950 700
rect 7600 650 8000 750
rect 7650 550 7750 650
rect 7850 550 7950 650
rect 7600 450 8000 550
rect -150 350 -50 450
rect 50 350 150 450
rect 250 350 350 400
rect 450 350 550 400
rect 650 350 750 400
rect 850 350 950 400
rect 1050 350 1150 400
rect 1250 350 1350 400
rect 1450 350 1550 400
rect 1650 350 1750 450
rect 3650 350 3750 450
rect 3850 350 3950 450
rect 4050 350 4150 450
rect 6050 350 6150 450
rect 6250 350 6350 400
rect 6450 350 6550 400
rect 6650 350 6750 400
rect 6850 350 6950 400
rect 7050 350 7150 400
rect 7250 350 7350 400
rect 7450 350 7550 400
rect 7650 350 7750 450
rect 7850 350 7950 450
rect -200 250 1800 350
rect 3600 250 4200 350
rect 6000 250 8000 350
rect -150 150 -50 250
rect 50 150 150 250
rect 250 150 350 250
rect 450 150 550 250
rect 650 150 750 250
rect 850 150 950 250
rect 1050 150 1150 250
rect 1250 150 1350 250
rect 1450 150 1550 250
rect 1650 150 1750 250
rect 1850 150 1950 200
rect 2050 150 2150 200
rect 2250 150 2350 200
rect 2450 150 2550 200
rect 2650 150 2750 200
rect 2850 150 2950 200
rect 3050 150 3150 200
rect 3250 150 3350 200
rect 3450 150 3550 200
rect 3650 150 3750 250
rect 3850 150 3950 250
rect 4050 150 4150 250
rect 4250 150 4350 200
rect 4450 150 4550 200
rect 4650 150 4750 200
rect 4850 150 4950 200
rect 5050 150 5150 200
rect 5250 150 5350 200
rect 5450 150 5550 200
rect 5650 150 5750 200
rect 5850 150 5950 200
rect 6050 150 6150 250
rect 6250 150 6350 250
rect 6450 150 6550 250
rect 6650 150 6750 250
rect 6850 150 6950 250
rect 7050 150 7150 250
rect 7250 150 7350 250
rect 7450 150 7550 250
rect 7650 150 7750 250
rect 7850 150 7950 250
rect -200 50 8000 150
rect -150 -50 -50 50
rect 50 -50 150 50
rect 250 -50 350 50
rect 450 -50 550 50
rect 650 -50 750 50
rect 850 -50 950 50
rect 1050 -50 1150 50
rect 1250 -50 1350 50
rect 1450 -50 1550 50
rect 1650 -50 1750 50
rect 1850 -50 1950 50
rect 2050 -50 2150 50
rect 2250 -50 2350 50
rect 2450 -50 2550 50
rect 2650 -50 2750 50
rect 2850 -50 2950 50
rect 3050 -50 3150 50
rect 3250 -50 3350 50
rect 3450 -50 3550 50
rect 3650 -50 3750 50
rect 3850 -50 3950 50
rect 4050 -50 4150 50
rect 4250 -50 4350 50
rect 4450 -50 4550 50
rect 4650 -50 4750 50
rect 4850 -50 4950 50
rect 5050 -50 5150 50
rect 5250 -50 5350 50
rect 5450 -50 5550 50
rect 5650 -50 5750 50
rect 5850 -50 5950 50
rect 6050 -50 6150 50
rect 6250 -50 6350 50
rect 6450 -50 6550 50
rect 6650 -50 6750 50
rect 6850 -50 6950 50
rect 7050 -50 7150 50
rect 7250 -50 7350 50
rect 7450 -50 7550 50
rect 7650 -50 7750 50
rect 7850 -50 7950 50
rect -200 -150 8000 -50
rect -150 -200 -50 -150
rect 50 -200 150 -150
rect 250 -200 350 -150
rect 450 -200 550 -150
rect 650 -200 750 -150
rect 850 -200 950 -150
rect 1050 -200 1150 -150
rect 1250 -200 1350 -150
rect 1450 -200 1550 -150
rect 1650 -200 1750 -150
rect 1850 -200 1950 -150
rect 2050 -200 2150 -150
rect 2250 -200 2350 -150
rect 2450 -200 2550 -150
rect 2650 -200 2750 -150
rect 2850 -200 2950 -150
rect 3050 -200 3150 -150
rect 3250 -200 3350 -150
rect 3450 -200 3550 -150
rect 3650 -200 3750 -150
rect 3850 -200 3950 -150
rect 4050 -200 4150 -150
rect 4250 -200 4350 -150
rect 4450 -200 4550 -150
rect 4650 -200 4750 -150
rect 4850 -200 4950 -150
rect 5050 -200 5150 -150
rect 5250 -200 5350 -150
rect 5450 -200 5550 -150
rect 5650 -200 5750 -150
rect 5850 -200 5950 -150
rect 6050 -200 6150 -150
rect 6250 -200 6350 -150
rect 6450 -200 6550 -150
rect 6650 -200 6750 -150
rect 6850 -200 6950 -150
rect 7050 -200 7150 -150
rect 7250 -200 7350 -150
rect 7450 -200 7550 -150
rect 7650 -200 7750 -150
rect 7850 -200 7950 -150
<< metal3 >>
rect 3250 3340 3350 3350
rect 3060 3260 3350 3340
rect 850 2340 950 2350
rect 850 2260 2140 2340
rect 850 2250 950 2260
rect 2060 2150 2140 2260
rect 1050 2140 1150 2150
rect 1050 2060 1740 2140
rect 1050 2050 1150 2060
rect 850 1850 950 1950
rect 850 1140 950 1150
rect 1060 1140 1140 2050
rect 1660 1350 1740 2060
rect 2050 2050 2150 2150
rect 3060 1750 3140 3260
rect 3250 3250 3350 3260
rect 4450 3340 4550 3350
rect 4450 3260 4740 3340
rect 4450 3250 4550 3260
rect 3250 3050 3350 3150
rect 4450 3050 4550 3150
rect 3050 1650 3150 1750
rect 1250 1340 1350 1350
rect 1650 1340 1750 1350
rect 1250 1260 1750 1340
rect 1250 1250 1350 1260
rect 1650 1250 1750 1260
rect 1660 1140 1740 1250
rect 3260 1140 3340 3050
rect 850 1060 3340 1140
rect 4460 1140 4540 3050
rect 4660 1750 4740 3260
rect 6850 2340 6950 2350
rect 5660 2260 6950 2340
rect 5660 2150 5740 2260
rect 6850 2250 6950 2260
rect 5650 2050 5750 2150
rect 6650 2140 6750 2150
rect 6060 2060 6750 2140
rect 4650 1650 4750 1750
rect 6060 1350 6140 2060
rect 6650 2050 6750 2060
rect 7050 2050 7150 2150
rect 6850 1850 6950 1950
rect 6050 1340 6150 1350
rect 6450 1340 6550 1350
rect 6050 1260 6550 1340
rect 6050 1250 6150 1260
rect 6450 1250 6550 1260
rect 6060 1140 6140 1250
rect 6850 1140 6950 1150
rect 4460 1060 6950 1140
rect 850 1050 950 1060
rect 1060 950 1140 1060
rect 2060 950 2140 1060
rect 5660 950 5740 1060
rect 6850 1050 6950 1060
rect 7060 950 7140 2050
rect 1050 940 1150 950
rect 1650 940 1750 950
rect 2050 940 2150 950
rect 3250 940 3350 950
rect 1050 860 2150 940
rect 1050 850 1150 860
rect 1650 850 1750 860
rect 1860 740 1940 860
rect 2050 850 2150 860
rect 3060 860 3350 940
rect 2060 750 2140 850
rect 2050 740 2150 750
rect 1860 660 2150 740
rect 2050 650 2150 660
rect 3060 540 3140 860
rect 3250 850 3350 860
rect 3450 940 3550 950
rect 4450 940 4550 950
rect 3450 860 4550 940
rect 3450 850 3550 860
rect 4450 850 4550 860
rect 5650 940 5750 950
rect 6050 940 6150 950
rect 6650 940 6750 950
rect 5650 860 6750 940
rect 5650 850 5750 860
rect 5660 750 5740 850
rect 3250 650 3350 750
rect 4450 650 4550 750
rect 5650 740 5750 750
rect 5860 740 5940 860
rect 6050 850 6150 860
rect 6650 850 6750 860
rect 7050 850 7150 950
rect 5650 660 5940 740
rect 5650 650 5750 660
rect 4460 540 4540 650
rect 3060 460 4540 540
<< metal4 >>
rect 860 1860 1140 1940
rect 1060 1340 1140 1860
rect 6660 1860 6940 1940
rect 6660 1340 6740 1860
rect 1060 1260 1340 1340
rect 1660 860 1740 1340
rect 3260 860 3540 940
rect 6060 860 6140 1340
rect 6460 1260 6740 1340
rect 3260 660 3340 860
use via_M1_M2_1_a  NoName_194 ~/A2G/A2G/magic/magic_layout/skywater130_microtemplates_dense
timestamp 1647525606
transform 1 0 3078 0 1 3364
box -32 -32 32 32
use via_M1_M2_1_b  NoName_195 ~/A2G/A2G/magic/magic_layout/skywater130_microtemplates_dense
timestamp 1647525606
transform 1 0 3078 0 1 3236
box -32 -32 32 32
use via_M1_M2_1_c  NoName_196 ~/A2G/A2G/magic/magic_layout/skywater130_microtemplates_dense
timestamp 1647525606
transform 1 0 3078 0 1 3492
box -32 -32 32 32
use via_M1_M2_1_d  NoName_197 ~/A2G/A2G/magic/magic_layout/skywater130_microtemplates_dense
timestamp 1647525606
transform 1 0 3078 0 1 3108
box -32 -32 32 32
use via_M1_M2_1_e  NoName_198 ~/A2G/A2G/magic/magic_layout/skywater130_microtemplates_dense
timestamp 1647525606
transform 1 0 4722 0 1 3364
box -32 -32 32 32
use via_M1_M2_1_f  NoName_199 ~/A2G/A2G/magic/magic_layout/skywater130_microtemplates_dense
timestamp 1647525606
transform 1 0 4722 0 1 3236
box -32 -32 32 32
use via_M1_M2_1_g  NoName_200 ~/A2G/A2G/magic/magic_layout/skywater130_microtemplates_dense
timestamp 1647525606
transform 1 0 4722 0 1 3492
box -32 -32 32 32
use via_M1_M2_1_h  NoName_201 ~/A2G/A2G/magic/magic_layout/skywater130_microtemplates_dense
timestamp 1647525606
transform 1 0 4722 0 1 3108
box -32 -32 32 32
use via_M1_M2_1_i  NoName_202 ~/A2G/A2G/magic/magic_layout/skywater130_microtemplates_dense
timestamp 1647525606
transform 1 0 1878 0 1 2100
box -32 -32 32 32
use via_M1_M2_1_j  NoName_203 ~/A2G/A2G/magic/magic_layout/skywater130_microtemplates_dense
timestamp 1647525606
transform 1 0 1878 0 1 2228
box -32 -32 32 32
use via_M1_M2_1_k  NoName_204 ~/A2G/A2G/magic/magic_layout/skywater130_microtemplates_dense
timestamp 1647525606
transform 1 0 1878 0 1 1972
box -32 -32 32 32
use via_M1_M2_1_l  NoName_205 ~/A2G/A2G/magic/magic_layout/skywater130_microtemplates_dense
timestamp 1647525606
transform 1 0 1878 0 1 2356
box -32 -32 32 32
use via_M1_M2_1_m  NoName_206 ~/A2G/A2G/magic/magic_layout/skywater130_microtemplates_dense
timestamp 1647525606
transform 1 0 1878 0 1 1844
box -32 -32 32 32
use via_M1_M2_1_n  NoName_207 ~/A2G/A2G/magic/magic_layout/skywater130_microtemplates_dense
timestamp 1647525606
transform 1 0 1878 0 1 2484
box -32 -32 32 32
use via_M1_M2_1_o  NoName_208 ~/A2G/A2G/magic/magic_layout/skywater130_microtemplates_dense
timestamp 1647525606
transform 1 0 1878 0 1 1716
box -32 -32 32 32
use via_M1_M2_1_p  NoName_209 ~/A2G/A2G/magic/magic_layout/skywater130_microtemplates_dense
timestamp 1647525606
transform 1 0 3522 0 1 2100
box -32 -32 32 32
use via_M1_M2_1_q  NoName_210 ~/A2G/A2G/magic/magic_layout/skywater130_microtemplates_dense
timestamp 1647525606
transform 1 0 3522 0 1 2228
box -32 -32 32 32
use via_M1_M2_1_r  NoName_211 ~/A2G/A2G/magic/magic_layout/skywater130_microtemplates_dense
timestamp 1647525606
transform 1 0 3522 0 1 1972
box -32 -32 32 32
use via_M1_M2_1_s  NoName_212 ~/A2G/A2G/magic/magic_layout/skywater130_microtemplates_dense
timestamp 1647525606
transform 1 0 3522 0 1 2356
box -32 -32 32 32
use via_M1_M2_1_t  NoName_213 ~/A2G/A2G/magic/magic_layout/skywater130_microtemplates_dense
timestamp 1647525606
transform 1 0 3522 0 1 1844
box -32 -32 32 32
use via_M1_M2_1_u  NoName_214 ~/A2G/A2G/magic/magic_layout/skywater130_microtemplates_dense
timestamp 1647525606
transform 1 0 3522 0 1 2484
box -32 -32 32 32
use via_M1_M2_1_v  NoName_215 ~/A2G/A2G/magic/magic_layout/skywater130_microtemplates_dense
timestamp 1647525606
transform 1 0 3522 0 1 1716
box -32 -32 32 32
use via_M1_M2_1_w  NoName_216 ~/A2G/A2G/magic/magic_layout/skywater130_microtemplates_dense
timestamp 1647525606
transform 1 0 4278 0 1 2100
box -32 -32 32 32
use via_M1_M2_1_x  NoName_217 ~/A2G/A2G/magic/magic_layout/skywater130_microtemplates_dense
timestamp 1647525606
transform 1 0 4278 0 1 2228
box -32 -32 32 32
use via_M1_M2_1_y  NoName_218 ~/A2G/A2G/magic/magic_layout/skywater130_microtemplates_dense
timestamp 1647525606
transform 1 0 4278 0 1 1972
box -32 -32 32 32
use via_M1_M2_1_z  NoName_219 ~/A2G/A2G/magic/magic_layout/skywater130_microtemplates_dense
timestamp 1647525606
transform 1 0 4278 0 1 2356
box -32 -32 32 32
use via_M1_M2_1_{  NoName_220 ~/A2G/A2G/magic/magic_layout/skywater130_microtemplates_dense
timestamp 1647525606
transform 1 0 4278 0 1 1844
box -32 -32 32 32
use via_M1_M2_1_|  NoName_221 ~/A2G/A2G/magic/magic_layout/skywater130_microtemplates_dense
timestamp 1647525606
transform 1 0 4278 0 1 2484
box -32 -32 32 32
use via_M1_M2_1_}  NoName_222 ~/A2G/A2G/magic/magic_layout/skywater130_microtemplates_dense
timestamp 1647525606
transform 1 0 4278 0 1 1716
box -32 -32 32 32
use via_M1_M2_1_~  NoName_223 ~/A2G/A2G/magic/magic_layout/skywater130_microtemplates_dense
timestamp 1647525606
transform 1 0 5922 0 1 2100
box -32 -32 32 32
use via_M1_M2_1_  NoName_224 ~/A2G/A2G/magic/magic_layout/skywater130_microtemplates_dense
timestamp 1647525606
transform 1 0 5922 0 1 2228
box -32 -32 32 32
use via_M1_M2_1_�  NoName_225 ~/A2G/A2G/magic/magic_layout/skywater130_microtemplates_dense
timestamp 1647525606
transform 1 0 5922 0 1 1972
box -32 -32 32 32
use via_M1_M2_1_�  NoName_226 ~/A2G/A2G/magic/magic_layout/skywater130_microtemplates_dense
timestamp 1647525606
transform 1 0 5922 0 1 2356
box -32 -32 32 32
use via_M1_M2_1_�  NoName_227 ~/A2G/A2G/magic/magic_layout/skywater130_microtemplates_dense
timestamp 1647525606
transform 1 0 5922 0 1 1844
box -32 -32 32 32
use via_M1_M2_1_�  NoName_228 ~/A2G/A2G/magic/magic_layout/skywater130_microtemplates_dense
timestamp 1647525606
transform 1 0 5922 0 1 2484
box -32 -32 32 32
use via_M1_M2_1_�  NoName_229 ~/A2G/A2G/magic/magic_layout/skywater130_microtemplates_dense
timestamp 1647525606
transform 1 0 5922 0 1 1716
box -32 -32 32 32
use via_M1_M2_1_�  NoName_230 ~/A2G/A2G/magic/magic_layout/skywater130_microtemplates_dense
timestamp 1647525606
transform 1 0 314 0 1 2164
box -32 -32 32 32
use via_M1_M2_1_�  NoName_231 ~/A2G/A2G/magic/magic_layout/skywater130_microtemplates_dense
timestamp 1647525606
transform 1 0 314 0 1 2036
box -32 -32 32 32
use via_M1_M2_1_�  NoName_232 ~/A2G/A2G/magic/magic_layout/skywater130_microtemplates_dense
timestamp 1647525606
transform 1 0 314 0 1 2292
box -32 -32 32 32
use via_M1_M2_1_�  NoName_233 ~/A2G/A2G/magic/magic_layout/skywater130_microtemplates_dense
timestamp 1647525606
transform 1 0 314 0 1 1906
box -32 -32 32 32
use via_M1_M2_1_�  NoName_234 ~/A2G/A2G/magic/magic_layout/skywater130_microtemplates_dense
timestamp 1647525606
transform 1 0 1486 0 1 2164
box -32 -32 32 32
use via_M1_M2_1_�  NoName_235 ~/A2G/A2G/magic/magic_layout/skywater130_microtemplates_dense
timestamp 1647525606
transform 1 0 1486 0 1 2036
box -32 -32 32 32
use via_M1_M2_1_�  NoName_236 ~/A2G/A2G/magic/magic_layout/skywater130_microtemplates_dense
timestamp 1647525606
transform 1 0 1486 0 1 2292
box -32 -32 32 32
use via_M1_M2_1_�  NoName_237 ~/A2G/A2G/magic/magic_layout/skywater130_microtemplates_dense
timestamp 1647525606
transform 1 0 1486 0 1 1906
box -32 -32 32 32
use via_M1_M2_1_�  NoName_238 ~/A2G/A2G/magic/magic_layout/skywater130_microtemplates_dense
timestamp 1647525606
transform 1 0 6314 0 1 2164
box -32 -32 32 32
use via_M1_M2_1_�  NoName_239 ~/A2G/A2G/magic/magic_layout/skywater130_microtemplates_dense
timestamp 1647525606
transform 1 0 6314 0 1 2036
box -32 -32 32 32
use via_M1_M2_1_�  NoName_240 ~/A2G/A2G/magic/magic_layout/skywater130_microtemplates_dense
timestamp 1647525606
transform 1 0 6314 0 1 2292
box -32 -32 32 32
use via_M1_M2_1_�  NoName_241 ~/A2G/A2G/magic/magic_layout/skywater130_microtemplates_dense
timestamp 1647525606
transform 1 0 6314 0 1 1906
box -32 -32 32 32
use via_M1_M2_1_�  NoName_242 ~/A2G/A2G/magic/magic_layout/skywater130_microtemplates_dense
timestamp 1647525606
transform 1 0 7486 0 1 2164
box -32 -32 32 32
use via_M1_M2_1_�  NoName_243 ~/A2G/A2G/magic/magic_layout/skywater130_microtemplates_dense
timestamp 1647525606
transform 1 0 7486 0 1 2036
box -32 -32 32 32
use via_M1_M2_1_�  NoName_244 ~/A2G/A2G/magic/magic_layout/skywater130_microtemplates_dense
timestamp 1647525606
transform 1 0 7486 0 1 2292
box -32 -32 32 32
use via_M1_M2_1_�  NoName_245 ~/A2G/A2G/magic/magic_layout/skywater130_microtemplates_dense
timestamp 1647525606
transform 1 0 7486 0 1 1906
box -32 -32 32 32
use via_M2_M3_0  NoName_246 ~/A2G/A2G/magic/magic_layout/skywater130_microtemplates_dense
timestamp 1647525786
transform 1 0 4500 0 1 3100
box -38 -38 38 38
use via_M2_M3_0  NoName_247
timestamp 1647525786
transform 1 0 6900 0 1 1100
box -38 -38 38 38
use via_M2_M3_0  NoName_250
timestamp 1647525786
transform 1 0 3300 0 1 3100
box -38 -38 38 38
use via_M2_M3_0  NoName_251
timestamp 1647525786
transform 1 0 900 0 1 1100
box -38 -38 38 38
use via_M2_M3_0  NoName_254
timestamp 1647525786
transform 1 0 2100 0 1 900
box -38 -38 38 38
use via_M2_M3_0  NoName_255
timestamp 1647525786
transform 1 0 900 0 1 1900
box -38 -38 38 38
use via_M3_M4_0  NoName_257 ~/A2G/A2G/magic/magic_layout/skywater130_microtemplates_dense
timestamp 1647526059
transform 1 0 1300 0 1 1300
box -38 -38 38 38
use via_M3_M4_0  NoName_258
timestamp 1647526059
transform 1 0 900 0 1 1900
box -38 -38 38 38
use via_M2_M3_0  NoName_260
timestamp 1647525786
transform 1 0 5700 0 1 900
box -38 -38 38 38
use via_M2_M3_0  NoName_261
timestamp 1647525786
transform 1 0 6900 0 1 1900
box -38 -38 38 38
use via_M3_M4_0  NoName_263
timestamp 1647526059
transform 1 0 6500 0 1 1300
box -38 -38 38 38
use via_M3_M4_0  NoName_264
timestamp 1647526059
transform 1 0 6900 0 1 1900
box -38 -38 38 38
use via_M2_M3_0  NoName_266
timestamp 1647525786
transform 1 0 5700 0 1 700
box -38 -38 38 38
use via_M2_M3_0  NoName_267
timestamp 1647525786
transform 1 0 6700 0 1 2100
box -38 -38 38 38
use via_M3_M4_0  NoName_269
timestamp 1647526059
transform 1 0 6100 0 1 900
box -38 -38 38 38
use via_M3_M4_0  NoName_270
timestamp 1647526059
transform 1 0 6100 0 1 1300
box -38 -38 38 38
use via_M2_M3_0  NoName_272
timestamp 1647525786
transform 1 0 2100 0 1 700
box -38 -38 38 38
use via_M2_M3_0  NoName_273
timestamp 1647525786
transform 1 0 1100 0 1 2100
box -38 -38 38 38
use via_M3_M4_0  NoName_275
timestamp 1647526059
transform 1 0 1700 0 1 900
box -38 -38 38 38
use via_M3_M4_0  NoName_276
timestamp 1647526059
transform 1 0 1700 0 1 1300
box -38 -38 38 38
use via_M2_M3_0  NoName_278
timestamp 1647525786
transform 1 0 1100 0 1 900
box -38 -38 38 38
use via_M2_M3_0  NoName_287
timestamp 1647525786
transform 1 0 6700 0 1 900
box -38 -38 38 38
use via_M2_M3_0  NoName_290
timestamp 1647525786
transform 1 0 3300 0 1 700
box -38 -38 38 38
use via_M2_M3_0  NoName_291
timestamp 1647525786
transform 1 0 4500 0 1 900
box -38 -38 38 38
use via_M3_M4_0  NoName_293
timestamp 1647526059
transform 1 0 3300 0 1 700
box -38 -38 38 38
use via_M3_M4_0  NoName_294
timestamp 1647526059
transform 1 0 3500 0 1 900
box -38 -38 38 38
use via_M2_M3_0  NoName_296
timestamp 1647525786
transform 1 0 4500 0 1 700
box -38 -38 38 38
use via_M2_M3_0  NoName_297
timestamp 1647525786
transform 1 0 3300 0 1 900
box -38 -38 38 38
use via_M2_M3_0  NoName_300
timestamp 1647525786
transform 1 0 4500 0 1 3300
box -38 -38 38 38
use via_M2_M3_0  NoName_301
timestamp 1647525786
transform 1 0 4700 0 1 1700
box -38 -38 38 38
use via_M2_M3_0  NoName_304
timestamp 1647525786
transform 1 0 3300 0 1 3300
box -38 -38 38 38
use via_M2_M3_0  NoName_305
timestamp 1647525786
transform 1 0 3100 0 1 1700
box -38 -38 38 38
use via_M2_M3_0  NoName_308
timestamp 1647525786
transform 1 0 2100 0 1 2100
box -38 -38 38 38
use via_M2_M3_0  NoName_309
timestamp 1647525786
transform 1 0 900 0 1 2300
box -38 -38 38 38
use via_M2_M3_0  NoName_312
timestamp 1647525786
transform 1 0 5700 0 1 2100
box -38 -38 38 38
use via_M2_M3_0  NoName_313
timestamp 1647525786
transform 1 0 6900 0 1 2300
box -38 -38 38 38
use via_M2_M3_0  NoName_316
timestamp 1647525786
transform 1 0 7100 0 1 900
box -38 -38 38 38
use via_M2_M3_0  NoName_317
timestamp 1647525786
transform 1 0 7100 0 1 2100
box -38 -38 38 38
use via_M1_M2_1  NoName_320 ~/A2G/A2G/magic/magic_layout/skywater130_microtemplates_dense
timestamp 1647525606
transform 1 0 4500 0 1 1150
box -32 -32 32 32
use via_M1_M2_1  NoName_321
timestamp 1647525606
transform 1 0 4700 0 1 1150
box -32 -32 32 32
use via_M1_M2_1  NoName_322
timestamp 1647525606
transform 1 0 4900 0 1 1150
box -32 -32 32 32
use via_M1_M2_1  NoName_323
timestamp 1647525606
transform 1 0 5100 0 1 1150
box -32 -32 32 32
use via_M1_M2_1  NoName_324
timestamp 1647525606
transform 1 0 5300 0 1 1150
box -32 -32 32 32
use via_M1_M2_1  NoName_325
timestamp 1647525606
transform 1 0 5500 0 1 1150
box -32 -32 32 32
use via_M1_M2_1  NoName_326
timestamp 1647525606
transform 1 0 5700 0 1 1150
box -32 -32 32 32
use via_M1_M2_1  NoName_327
timestamp 1647525606
transform 1 0 2100 0 1 1150
box -32 -32 32 32
use via_M1_M2_1  NoName_328
timestamp 1647525606
transform 1 0 2300 0 1 1150
box -32 -32 32 32
use via_M1_M2_1  NoName_329
timestamp 1647525606
transform 1 0 2500 0 1 1150
box -32 -32 32 32
use via_M1_M2_1  NoName_330
timestamp 1647525606
transform 1 0 2700 0 1 1150
box -32 -32 32 32
use via_M1_M2_1  NoName_331
timestamp 1647525606
transform 1 0 2900 0 1 1150
box -32 -32 32 32
use via_M1_M2_1  NoName_332
timestamp 1647525606
transform 1 0 3100 0 1 1150
box -32 -32 32 32
use via_M1_M2_1  NoName_333
timestamp 1647525606
transform 1 0 3300 0 1 1150
box -32 -32 32 32
use via_M1_M2_1  NoName_334
timestamp 1647525606
transform 1 0 6900 0 1 550
box -32 -32 32 32
use via_M1_M2_1  NoName_335
timestamp 1647525606
transform 1 0 900 0 1 550
box -32 -32 32 32
use XM2  XM2 ~/A2G/A2G/magic/magic_layout/pcell
timestamp 1686266349
transform 1 0 900 0 1 900
box -639 -364 639 364
use XM3  XM3 ~/A2G/A2G/magic/magic_layout/pcell
timestamp 1686266349
transform 1 0 6900 0 1 900
box -639 -364 639 364
use XMdiff  XMdiff ~/A2G/A2G/magic/magic_layout/pcell
timestamp 1686266346
transform -1 0 3900 0 -1 3300
box -875 -359 875 359
use XMinn  XMinn ~/A2G/A2G/magic/magic_layout/pcell
timestamp 1686266346
transform 1 0 2700 0 1 2100
box -875 -539 875 539
use XMinp  XMinp ~/A2G/A2G/magic/magic_layout/pcell
timestamp 1686266347
transform 1 0 5100 0 1 2100
box -875 -539 875 539
use XMl1  XMl1 ~/A2G/A2G/magic/magic_layout/pcell
timestamp 1686266350
transform -1 0 900 0 -1 2100
box -639 -359 639 359
use XMl2  XMl2 ~/A2G/A2G/magic/magic_layout/pcell
timestamp 1686266350
transform -1 0 6900 0 -1 2100
box -639 -359 639 359
use XMl3  XMl3 ~/A2G/A2G/magic/magic_layout/pcell
timestamp 1686266348
transform -1 0 2700 0 -1 700
box -875 -364 875 364
use XMl4  XMl4 ~/A2G/A2G/magic/magic_layout/pcell
timestamp 1686266348
transform -1 0 5100 0 -1 700
box -875 -364 875 364
<< labels >>
flabel metal3 3100 1100 3100 1100 0 FreeSans 1600 0 0 0 clk
flabel metal3 7100 1500 7100 1500 0 FreeSans 1600 0 0 0 outp
flabel metal3 3700 900 3700 900 0 FreeSans 1600 0 0 0 outn
flabel metal2 2700 2500 2700 2500 0 FreeSans 1600 0 0 0 vn
flabel metal2 5100 2500 5100 2500 0 FreeSans 1600 0 0 0 vp
flabel metal1 5100 500 5100 500 0 FreeSans 1600 0 0 0 vdd
flabel metal1 2700 500 2700 500 0 FreeSans 1600 0 0 0 vdd
flabel metal2 6900 700 6900 700 0 FreeSans 1600 0 0 0 vdd
flabel metal2 900 700 900 700 0 FreeSans 1600 0 0 0 vdd
flabel metal2 3900 3500 3900 3500 0 FreeSans 1600 0 0 0 vss
<< end >>
