magic
tech sky130A
timestamp 1680002671
<< error_p >>
rect -19 14 19 19
rect -19 -14 -14 14
rect -19 -19 19 -14
<< metal2 >>
rect -19 14 19 19
rect -19 -14 -14 14
rect 14 -14 19 14
rect -19 -19 19 -14
<< via2 >>
rect -14 -14 14 14
<< metal3 >>
rect -19 14 19 19
rect -19 -14 -14 14
rect 14 -14 19 14
rect -19 -19 19 -14
<< end >>
