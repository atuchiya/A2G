magic
tech sky130A
magscale 1 2
timestamp 1680002671
<< error_p >>
rect -991 391 -929 397
rect -863 391 -801 397
rect -735 391 -673 397
rect -607 391 -545 397
rect -479 391 -417 397
rect -351 391 -289 397
rect -223 391 -161 397
rect -95 391 -33 397
rect 33 391 95 397
rect 161 391 223 397
rect 289 391 351 397
rect 417 391 479 397
rect 545 391 607 397
rect 673 391 735 397
rect 801 391 863 397
rect 929 391 991 397
rect -991 357 -977 391
rect -863 357 -849 391
rect -735 357 -721 391
rect -607 357 -593 391
rect -479 357 -465 391
rect -351 357 -337 391
rect -223 357 -209 391
rect -95 357 -81 391
rect 33 357 47 391
rect 161 357 175 391
rect 289 357 303 391
rect 417 357 431 391
rect 545 357 559 391
rect 673 357 687 391
rect 801 357 815 391
rect 929 357 943 391
rect -991 351 -929 357
rect -863 351 -801 357
rect -735 351 -673 357
rect -607 351 -545 357
rect -479 351 -417 357
rect -351 351 -289 357
rect -223 351 -161 357
rect -95 351 -33 357
rect 33 351 95 357
rect 161 351 223 357
rect 289 351 351 357
rect 417 351 479 357
rect 545 351 607 357
rect 673 351 735 357
rect 801 351 863 357
rect 929 351 991 357
<< pwell >>
rect -1181 -519 1181 519
<< nmoslvt >>
rect -995 -381 -925 319
rect -867 -381 -797 319
rect -739 -381 -669 319
rect -611 -381 -541 319
rect -483 -381 -413 319
rect -355 -381 -285 319
rect -227 -381 -157 319
rect -99 -381 -29 319
rect 29 -381 99 319
rect 157 -381 227 319
rect 285 -381 355 319
rect 413 -381 483 319
rect 541 -381 611 319
rect 669 -381 739 319
rect 797 -381 867 319
rect 925 -381 995 319
<< ndiff >>
rect -1053 292 -995 319
rect -1053 258 -1041 292
rect -1007 258 -995 292
rect -1053 224 -995 258
rect -1053 190 -1041 224
rect -1007 190 -995 224
rect -1053 156 -995 190
rect -1053 122 -1041 156
rect -1007 122 -995 156
rect -1053 88 -995 122
rect -1053 54 -1041 88
rect -1007 54 -995 88
rect -1053 20 -995 54
rect -1053 -14 -1041 20
rect -1007 -14 -995 20
rect -1053 -48 -995 -14
rect -1053 -82 -1041 -48
rect -1007 -82 -995 -48
rect -1053 -116 -995 -82
rect -1053 -150 -1041 -116
rect -1007 -150 -995 -116
rect -1053 -184 -995 -150
rect -1053 -218 -1041 -184
rect -1007 -218 -995 -184
rect -1053 -252 -995 -218
rect -1053 -286 -1041 -252
rect -1007 -286 -995 -252
rect -1053 -320 -995 -286
rect -1053 -354 -1041 -320
rect -1007 -354 -995 -320
rect -1053 -381 -995 -354
rect -925 292 -867 319
rect -925 258 -913 292
rect -879 258 -867 292
rect -925 224 -867 258
rect -925 190 -913 224
rect -879 190 -867 224
rect -925 156 -867 190
rect -925 122 -913 156
rect -879 122 -867 156
rect -925 88 -867 122
rect -925 54 -913 88
rect -879 54 -867 88
rect -925 20 -867 54
rect -925 -14 -913 20
rect -879 -14 -867 20
rect -925 -48 -867 -14
rect -925 -82 -913 -48
rect -879 -82 -867 -48
rect -925 -116 -867 -82
rect -925 -150 -913 -116
rect -879 -150 -867 -116
rect -925 -184 -867 -150
rect -925 -218 -913 -184
rect -879 -218 -867 -184
rect -925 -252 -867 -218
rect -925 -286 -913 -252
rect -879 -286 -867 -252
rect -925 -320 -867 -286
rect -925 -354 -913 -320
rect -879 -354 -867 -320
rect -925 -381 -867 -354
rect -797 292 -739 319
rect -797 258 -785 292
rect -751 258 -739 292
rect -797 224 -739 258
rect -797 190 -785 224
rect -751 190 -739 224
rect -797 156 -739 190
rect -797 122 -785 156
rect -751 122 -739 156
rect -797 88 -739 122
rect -797 54 -785 88
rect -751 54 -739 88
rect -797 20 -739 54
rect -797 -14 -785 20
rect -751 -14 -739 20
rect -797 -48 -739 -14
rect -797 -82 -785 -48
rect -751 -82 -739 -48
rect -797 -116 -739 -82
rect -797 -150 -785 -116
rect -751 -150 -739 -116
rect -797 -184 -739 -150
rect -797 -218 -785 -184
rect -751 -218 -739 -184
rect -797 -252 -739 -218
rect -797 -286 -785 -252
rect -751 -286 -739 -252
rect -797 -320 -739 -286
rect -797 -354 -785 -320
rect -751 -354 -739 -320
rect -797 -381 -739 -354
rect -669 292 -611 319
rect -669 258 -657 292
rect -623 258 -611 292
rect -669 224 -611 258
rect -669 190 -657 224
rect -623 190 -611 224
rect -669 156 -611 190
rect -669 122 -657 156
rect -623 122 -611 156
rect -669 88 -611 122
rect -669 54 -657 88
rect -623 54 -611 88
rect -669 20 -611 54
rect -669 -14 -657 20
rect -623 -14 -611 20
rect -669 -48 -611 -14
rect -669 -82 -657 -48
rect -623 -82 -611 -48
rect -669 -116 -611 -82
rect -669 -150 -657 -116
rect -623 -150 -611 -116
rect -669 -184 -611 -150
rect -669 -218 -657 -184
rect -623 -218 -611 -184
rect -669 -252 -611 -218
rect -669 -286 -657 -252
rect -623 -286 -611 -252
rect -669 -320 -611 -286
rect -669 -354 -657 -320
rect -623 -354 -611 -320
rect -669 -381 -611 -354
rect -541 292 -483 319
rect -541 258 -529 292
rect -495 258 -483 292
rect -541 224 -483 258
rect -541 190 -529 224
rect -495 190 -483 224
rect -541 156 -483 190
rect -541 122 -529 156
rect -495 122 -483 156
rect -541 88 -483 122
rect -541 54 -529 88
rect -495 54 -483 88
rect -541 20 -483 54
rect -541 -14 -529 20
rect -495 -14 -483 20
rect -541 -48 -483 -14
rect -541 -82 -529 -48
rect -495 -82 -483 -48
rect -541 -116 -483 -82
rect -541 -150 -529 -116
rect -495 -150 -483 -116
rect -541 -184 -483 -150
rect -541 -218 -529 -184
rect -495 -218 -483 -184
rect -541 -252 -483 -218
rect -541 -286 -529 -252
rect -495 -286 -483 -252
rect -541 -320 -483 -286
rect -541 -354 -529 -320
rect -495 -354 -483 -320
rect -541 -381 -483 -354
rect -413 292 -355 319
rect -413 258 -401 292
rect -367 258 -355 292
rect -413 224 -355 258
rect -413 190 -401 224
rect -367 190 -355 224
rect -413 156 -355 190
rect -413 122 -401 156
rect -367 122 -355 156
rect -413 88 -355 122
rect -413 54 -401 88
rect -367 54 -355 88
rect -413 20 -355 54
rect -413 -14 -401 20
rect -367 -14 -355 20
rect -413 -48 -355 -14
rect -413 -82 -401 -48
rect -367 -82 -355 -48
rect -413 -116 -355 -82
rect -413 -150 -401 -116
rect -367 -150 -355 -116
rect -413 -184 -355 -150
rect -413 -218 -401 -184
rect -367 -218 -355 -184
rect -413 -252 -355 -218
rect -413 -286 -401 -252
rect -367 -286 -355 -252
rect -413 -320 -355 -286
rect -413 -354 -401 -320
rect -367 -354 -355 -320
rect -413 -381 -355 -354
rect -285 292 -227 319
rect -285 258 -273 292
rect -239 258 -227 292
rect -285 224 -227 258
rect -285 190 -273 224
rect -239 190 -227 224
rect -285 156 -227 190
rect -285 122 -273 156
rect -239 122 -227 156
rect -285 88 -227 122
rect -285 54 -273 88
rect -239 54 -227 88
rect -285 20 -227 54
rect -285 -14 -273 20
rect -239 -14 -227 20
rect -285 -48 -227 -14
rect -285 -82 -273 -48
rect -239 -82 -227 -48
rect -285 -116 -227 -82
rect -285 -150 -273 -116
rect -239 -150 -227 -116
rect -285 -184 -227 -150
rect -285 -218 -273 -184
rect -239 -218 -227 -184
rect -285 -252 -227 -218
rect -285 -286 -273 -252
rect -239 -286 -227 -252
rect -285 -320 -227 -286
rect -285 -354 -273 -320
rect -239 -354 -227 -320
rect -285 -381 -227 -354
rect -157 292 -99 319
rect -157 258 -145 292
rect -111 258 -99 292
rect -157 224 -99 258
rect -157 190 -145 224
rect -111 190 -99 224
rect -157 156 -99 190
rect -157 122 -145 156
rect -111 122 -99 156
rect -157 88 -99 122
rect -157 54 -145 88
rect -111 54 -99 88
rect -157 20 -99 54
rect -157 -14 -145 20
rect -111 -14 -99 20
rect -157 -48 -99 -14
rect -157 -82 -145 -48
rect -111 -82 -99 -48
rect -157 -116 -99 -82
rect -157 -150 -145 -116
rect -111 -150 -99 -116
rect -157 -184 -99 -150
rect -157 -218 -145 -184
rect -111 -218 -99 -184
rect -157 -252 -99 -218
rect -157 -286 -145 -252
rect -111 -286 -99 -252
rect -157 -320 -99 -286
rect -157 -354 -145 -320
rect -111 -354 -99 -320
rect -157 -381 -99 -354
rect -29 292 29 319
rect -29 258 -17 292
rect 17 258 29 292
rect -29 224 29 258
rect -29 190 -17 224
rect 17 190 29 224
rect -29 156 29 190
rect -29 122 -17 156
rect 17 122 29 156
rect -29 88 29 122
rect -29 54 -17 88
rect 17 54 29 88
rect -29 20 29 54
rect -29 -14 -17 20
rect 17 -14 29 20
rect -29 -48 29 -14
rect -29 -82 -17 -48
rect 17 -82 29 -48
rect -29 -116 29 -82
rect -29 -150 -17 -116
rect 17 -150 29 -116
rect -29 -184 29 -150
rect -29 -218 -17 -184
rect 17 -218 29 -184
rect -29 -252 29 -218
rect -29 -286 -17 -252
rect 17 -286 29 -252
rect -29 -320 29 -286
rect -29 -354 -17 -320
rect 17 -354 29 -320
rect -29 -381 29 -354
rect 99 292 157 319
rect 99 258 111 292
rect 145 258 157 292
rect 99 224 157 258
rect 99 190 111 224
rect 145 190 157 224
rect 99 156 157 190
rect 99 122 111 156
rect 145 122 157 156
rect 99 88 157 122
rect 99 54 111 88
rect 145 54 157 88
rect 99 20 157 54
rect 99 -14 111 20
rect 145 -14 157 20
rect 99 -48 157 -14
rect 99 -82 111 -48
rect 145 -82 157 -48
rect 99 -116 157 -82
rect 99 -150 111 -116
rect 145 -150 157 -116
rect 99 -184 157 -150
rect 99 -218 111 -184
rect 145 -218 157 -184
rect 99 -252 157 -218
rect 99 -286 111 -252
rect 145 -286 157 -252
rect 99 -320 157 -286
rect 99 -354 111 -320
rect 145 -354 157 -320
rect 99 -381 157 -354
rect 227 292 285 319
rect 227 258 239 292
rect 273 258 285 292
rect 227 224 285 258
rect 227 190 239 224
rect 273 190 285 224
rect 227 156 285 190
rect 227 122 239 156
rect 273 122 285 156
rect 227 88 285 122
rect 227 54 239 88
rect 273 54 285 88
rect 227 20 285 54
rect 227 -14 239 20
rect 273 -14 285 20
rect 227 -48 285 -14
rect 227 -82 239 -48
rect 273 -82 285 -48
rect 227 -116 285 -82
rect 227 -150 239 -116
rect 273 -150 285 -116
rect 227 -184 285 -150
rect 227 -218 239 -184
rect 273 -218 285 -184
rect 227 -252 285 -218
rect 227 -286 239 -252
rect 273 -286 285 -252
rect 227 -320 285 -286
rect 227 -354 239 -320
rect 273 -354 285 -320
rect 227 -381 285 -354
rect 355 292 413 319
rect 355 258 367 292
rect 401 258 413 292
rect 355 224 413 258
rect 355 190 367 224
rect 401 190 413 224
rect 355 156 413 190
rect 355 122 367 156
rect 401 122 413 156
rect 355 88 413 122
rect 355 54 367 88
rect 401 54 413 88
rect 355 20 413 54
rect 355 -14 367 20
rect 401 -14 413 20
rect 355 -48 413 -14
rect 355 -82 367 -48
rect 401 -82 413 -48
rect 355 -116 413 -82
rect 355 -150 367 -116
rect 401 -150 413 -116
rect 355 -184 413 -150
rect 355 -218 367 -184
rect 401 -218 413 -184
rect 355 -252 413 -218
rect 355 -286 367 -252
rect 401 -286 413 -252
rect 355 -320 413 -286
rect 355 -354 367 -320
rect 401 -354 413 -320
rect 355 -381 413 -354
rect 483 292 541 319
rect 483 258 495 292
rect 529 258 541 292
rect 483 224 541 258
rect 483 190 495 224
rect 529 190 541 224
rect 483 156 541 190
rect 483 122 495 156
rect 529 122 541 156
rect 483 88 541 122
rect 483 54 495 88
rect 529 54 541 88
rect 483 20 541 54
rect 483 -14 495 20
rect 529 -14 541 20
rect 483 -48 541 -14
rect 483 -82 495 -48
rect 529 -82 541 -48
rect 483 -116 541 -82
rect 483 -150 495 -116
rect 529 -150 541 -116
rect 483 -184 541 -150
rect 483 -218 495 -184
rect 529 -218 541 -184
rect 483 -252 541 -218
rect 483 -286 495 -252
rect 529 -286 541 -252
rect 483 -320 541 -286
rect 483 -354 495 -320
rect 529 -354 541 -320
rect 483 -381 541 -354
rect 611 292 669 319
rect 611 258 623 292
rect 657 258 669 292
rect 611 224 669 258
rect 611 190 623 224
rect 657 190 669 224
rect 611 156 669 190
rect 611 122 623 156
rect 657 122 669 156
rect 611 88 669 122
rect 611 54 623 88
rect 657 54 669 88
rect 611 20 669 54
rect 611 -14 623 20
rect 657 -14 669 20
rect 611 -48 669 -14
rect 611 -82 623 -48
rect 657 -82 669 -48
rect 611 -116 669 -82
rect 611 -150 623 -116
rect 657 -150 669 -116
rect 611 -184 669 -150
rect 611 -218 623 -184
rect 657 -218 669 -184
rect 611 -252 669 -218
rect 611 -286 623 -252
rect 657 -286 669 -252
rect 611 -320 669 -286
rect 611 -354 623 -320
rect 657 -354 669 -320
rect 611 -381 669 -354
rect 739 292 797 319
rect 739 258 751 292
rect 785 258 797 292
rect 739 224 797 258
rect 739 190 751 224
rect 785 190 797 224
rect 739 156 797 190
rect 739 122 751 156
rect 785 122 797 156
rect 739 88 797 122
rect 739 54 751 88
rect 785 54 797 88
rect 739 20 797 54
rect 739 -14 751 20
rect 785 -14 797 20
rect 739 -48 797 -14
rect 739 -82 751 -48
rect 785 -82 797 -48
rect 739 -116 797 -82
rect 739 -150 751 -116
rect 785 -150 797 -116
rect 739 -184 797 -150
rect 739 -218 751 -184
rect 785 -218 797 -184
rect 739 -252 797 -218
rect 739 -286 751 -252
rect 785 -286 797 -252
rect 739 -320 797 -286
rect 739 -354 751 -320
rect 785 -354 797 -320
rect 739 -381 797 -354
rect 867 292 925 319
rect 867 258 879 292
rect 913 258 925 292
rect 867 224 925 258
rect 867 190 879 224
rect 913 190 925 224
rect 867 156 925 190
rect 867 122 879 156
rect 913 122 925 156
rect 867 88 925 122
rect 867 54 879 88
rect 913 54 925 88
rect 867 20 925 54
rect 867 -14 879 20
rect 913 -14 925 20
rect 867 -48 925 -14
rect 867 -82 879 -48
rect 913 -82 925 -48
rect 867 -116 925 -82
rect 867 -150 879 -116
rect 913 -150 925 -116
rect 867 -184 925 -150
rect 867 -218 879 -184
rect 913 -218 925 -184
rect 867 -252 925 -218
rect 867 -286 879 -252
rect 913 -286 925 -252
rect 867 -320 925 -286
rect 867 -354 879 -320
rect 913 -354 925 -320
rect 867 -381 925 -354
rect 995 292 1053 319
rect 995 258 1007 292
rect 1041 258 1053 292
rect 995 224 1053 258
rect 995 190 1007 224
rect 1041 190 1053 224
rect 995 156 1053 190
rect 995 122 1007 156
rect 1041 122 1053 156
rect 995 88 1053 122
rect 995 54 1007 88
rect 1041 54 1053 88
rect 995 20 1053 54
rect 995 -14 1007 20
rect 1041 -14 1053 20
rect 995 -48 1053 -14
rect 995 -82 1007 -48
rect 1041 -82 1053 -48
rect 995 -116 1053 -82
rect 995 -150 1007 -116
rect 1041 -150 1053 -116
rect 995 -184 1053 -150
rect 995 -218 1007 -184
rect 1041 -218 1053 -184
rect 995 -252 1053 -218
rect 995 -286 1007 -252
rect 1041 -286 1053 -252
rect 995 -320 1053 -286
rect 995 -354 1007 -320
rect 1041 -354 1053 -320
rect 995 -381 1053 -354
<< ndiffc >>
rect -1041 258 -1007 292
rect -1041 190 -1007 224
rect -1041 122 -1007 156
rect -1041 54 -1007 88
rect -1041 -14 -1007 20
rect -1041 -82 -1007 -48
rect -1041 -150 -1007 -116
rect -1041 -218 -1007 -184
rect -1041 -286 -1007 -252
rect -1041 -354 -1007 -320
rect -913 258 -879 292
rect -913 190 -879 224
rect -913 122 -879 156
rect -913 54 -879 88
rect -913 -14 -879 20
rect -913 -82 -879 -48
rect -913 -150 -879 -116
rect -913 -218 -879 -184
rect -913 -286 -879 -252
rect -913 -354 -879 -320
rect -785 258 -751 292
rect -785 190 -751 224
rect -785 122 -751 156
rect -785 54 -751 88
rect -785 -14 -751 20
rect -785 -82 -751 -48
rect -785 -150 -751 -116
rect -785 -218 -751 -184
rect -785 -286 -751 -252
rect -785 -354 -751 -320
rect -657 258 -623 292
rect -657 190 -623 224
rect -657 122 -623 156
rect -657 54 -623 88
rect -657 -14 -623 20
rect -657 -82 -623 -48
rect -657 -150 -623 -116
rect -657 -218 -623 -184
rect -657 -286 -623 -252
rect -657 -354 -623 -320
rect -529 258 -495 292
rect -529 190 -495 224
rect -529 122 -495 156
rect -529 54 -495 88
rect -529 -14 -495 20
rect -529 -82 -495 -48
rect -529 -150 -495 -116
rect -529 -218 -495 -184
rect -529 -286 -495 -252
rect -529 -354 -495 -320
rect -401 258 -367 292
rect -401 190 -367 224
rect -401 122 -367 156
rect -401 54 -367 88
rect -401 -14 -367 20
rect -401 -82 -367 -48
rect -401 -150 -367 -116
rect -401 -218 -367 -184
rect -401 -286 -367 -252
rect -401 -354 -367 -320
rect -273 258 -239 292
rect -273 190 -239 224
rect -273 122 -239 156
rect -273 54 -239 88
rect -273 -14 -239 20
rect -273 -82 -239 -48
rect -273 -150 -239 -116
rect -273 -218 -239 -184
rect -273 -286 -239 -252
rect -273 -354 -239 -320
rect -145 258 -111 292
rect -145 190 -111 224
rect -145 122 -111 156
rect -145 54 -111 88
rect -145 -14 -111 20
rect -145 -82 -111 -48
rect -145 -150 -111 -116
rect -145 -218 -111 -184
rect -145 -286 -111 -252
rect -145 -354 -111 -320
rect -17 258 17 292
rect -17 190 17 224
rect -17 122 17 156
rect -17 54 17 88
rect -17 -14 17 20
rect -17 -82 17 -48
rect -17 -150 17 -116
rect -17 -218 17 -184
rect -17 -286 17 -252
rect -17 -354 17 -320
rect 111 258 145 292
rect 111 190 145 224
rect 111 122 145 156
rect 111 54 145 88
rect 111 -14 145 20
rect 111 -82 145 -48
rect 111 -150 145 -116
rect 111 -218 145 -184
rect 111 -286 145 -252
rect 111 -354 145 -320
rect 239 258 273 292
rect 239 190 273 224
rect 239 122 273 156
rect 239 54 273 88
rect 239 -14 273 20
rect 239 -82 273 -48
rect 239 -150 273 -116
rect 239 -218 273 -184
rect 239 -286 273 -252
rect 239 -354 273 -320
rect 367 258 401 292
rect 367 190 401 224
rect 367 122 401 156
rect 367 54 401 88
rect 367 -14 401 20
rect 367 -82 401 -48
rect 367 -150 401 -116
rect 367 -218 401 -184
rect 367 -286 401 -252
rect 367 -354 401 -320
rect 495 258 529 292
rect 495 190 529 224
rect 495 122 529 156
rect 495 54 529 88
rect 495 -14 529 20
rect 495 -82 529 -48
rect 495 -150 529 -116
rect 495 -218 529 -184
rect 495 -286 529 -252
rect 495 -354 529 -320
rect 623 258 657 292
rect 623 190 657 224
rect 623 122 657 156
rect 623 54 657 88
rect 623 -14 657 20
rect 623 -82 657 -48
rect 623 -150 657 -116
rect 623 -218 657 -184
rect 623 -286 657 -252
rect 623 -354 657 -320
rect 751 258 785 292
rect 751 190 785 224
rect 751 122 785 156
rect 751 54 785 88
rect 751 -14 785 20
rect 751 -82 785 -48
rect 751 -150 785 -116
rect 751 -218 785 -184
rect 751 -286 785 -252
rect 751 -354 785 -320
rect 879 258 913 292
rect 879 190 913 224
rect 879 122 913 156
rect 879 54 913 88
rect 879 -14 913 20
rect 879 -82 913 -48
rect 879 -150 913 -116
rect 879 -218 913 -184
rect 879 -286 913 -252
rect 879 -354 913 -320
rect 1007 258 1041 292
rect 1007 190 1041 224
rect 1007 122 1041 156
rect 1007 54 1041 88
rect 1007 -14 1041 20
rect 1007 -82 1041 -48
rect 1007 -150 1041 -116
rect 1007 -218 1041 -184
rect 1007 -286 1041 -252
rect 1007 -354 1041 -320
<< psubdiff >>
rect -1155 459 -1037 493
rect -1003 459 -969 493
rect -935 459 -901 493
rect -867 459 -833 493
rect -799 459 -765 493
rect -731 459 -697 493
rect -663 459 -629 493
rect -595 459 -561 493
rect -527 459 -493 493
rect -459 459 -425 493
rect -391 459 -357 493
rect -323 459 -289 493
rect -255 459 -221 493
rect -187 459 -153 493
rect -119 459 -85 493
rect -51 459 -17 493
rect 17 459 51 493
rect 85 459 119 493
rect 153 459 187 493
rect 221 459 255 493
rect 289 459 323 493
rect 357 459 391 493
rect 425 459 459 493
rect 493 459 527 493
rect 561 459 595 493
rect 629 459 663 493
rect 697 459 731 493
rect 765 459 799 493
rect 833 459 867 493
rect 901 459 935 493
rect 969 459 1003 493
rect 1037 459 1155 493
rect -1155 391 -1121 459
rect -1155 323 -1121 357
rect 1121 391 1155 459
rect 1121 323 1155 357
rect -1155 255 -1121 289
rect -1155 187 -1121 221
rect -1155 119 -1121 153
rect -1155 51 -1121 85
rect -1155 -17 -1121 17
rect -1155 -85 -1121 -51
rect -1155 -153 -1121 -119
rect -1155 -221 -1121 -187
rect -1155 -289 -1121 -255
rect -1155 -357 -1121 -323
rect 1121 255 1155 289
rect 1121 187 1155 221
rect 1121 119 1155 153
rect 1121 51 1155 85
rect 1121 -17 1155 17
rect 1121 -85 1155 -51
rect 1121 -153 1155 -119
rect 1121 -221 1155 -187
rect 1121 -289 1155 -255
rect 1121 -357 1155 -323
rect -1155 -459 -1121 -391
rect 1121 -459 1155 -391
rect -1155 -493 -1037 -459
rect -1003 -493 -969 -459
rect -935 -493 -901 -459
rect -867 -493 -833 -459
rect -799 -493 -765 -459
rect -731 -493 -697 -459
rect -663 -493 -629 -459
rect -595 -493 -561 -459
rect -527 -493 -493 -459
rect -459 -493 -425 -459
rect -391 -493 -357 -459
rect -323 -493 -289 -459
rect -255 -493 -221 -459
rect -187 -493 -153 -459
rect -119 -493 -85 -459
rect -51 -493 -17 -459
rect 17 -493 51 -459
rect 85 -493 119 -459
rect 153 -493 187 -459
rect 221 -493 255 -459
rect 289 -493 323 -459
rect 357 -493 391 -459
rect 425 -493 459 -459
rect 493 -493 527 -459
rect 561 -493 595 -459
rect 629 -493 663 -459
rect 697 -493 731 -459
rect 765 -493 799 -459
rect 833 -493 867 -459
rect 901 -493 935 -459
rect 969 -493 1003 -459
rect 1037 -493 1155 -459
<< psubdiffcont >>
rect -1037 459 -1003 493
rect -969 459 -935 493
rect -901 459 -867 493
rect -833 459 -799 493
rect -765 459 -731 493
rect -697 459 -663 493
rect -629 459 -595 493
rect -561 459 -527 493
rect -493 459 -459 493
rect -425 459 -391 493
rect -357 459 -323 493
rect -289 459 -255 493
rect -221 459 -187 493
rect -153 459 -119 493
rect -85 459 -51 493
rect -17 459 17 493
rect 51 459 85 493
rect 119 459 153 493
rect 187 459 221 493
rect 255 459 289 493
rect 323 459 357 493
rect 391 459 425 493
rect 459 459 493 493
rect 527 459 561 493
rect 595 459 629 493
rect 663 459 697 493
rect 731 459 765 493
rect 799 459 833 493
rect 867 459 901 493
rect 935 459 969 493
rect 1003 459 1037 493
rect -1155 357 -1121 391
rect -1155 289 -1121 323
rect 1121 357 1155 391
rect -1155 221 -1121 255
rect -1155 153 -1121 187
rect -1155 85 -1121 119
rect -1155 17 -1121 51
rect -1155 -51 -1121 -17
rect -1155 -119 -1121 -85
rect -1155 -187 -1121 -153
rect -1155 -255 -1121 -221
rect -1155 -323 -1121 -289
rect -1155 -391 -1121 -357
rect 1121 289 1155 323
rect 1121 221 1155 255
rect 1121 153 1155 187
rect 1121 85 1155 119
rect 1121 17 1155 51
rect 1121 -51 1155 -17
rect 1121 -119 1155 -85
rect 1121 -187 1155 -153
rect 1121 -255 1155 -221
rect 1121 -323 1155 -289
rect 1121 -391 1155 -357
rect -1037 -493 -1003 -459
rect -969 -493 -935 -459
rect -901 -493 -867 -459
rect -833 -493 -799 -459
rect -765 -493 -731 -459
rect -697 -493 -663 -459
rect -629 -493 -595 -459
rect -561 -493 -527 -459
rect -493 -493 -459 -459
rect -425 -493 -391 -459
rect -357 -493 -323 -459
rect -289 -493 -255 -459
rect -221 -493 -187 -459
rect -153 -493 -119 -459
rect -85 -493 -51 -459
rect -17 -493 17 -459
rect 51 -493 85 -459
rect 119 -493 153 -459
rect 187 -493 221 -459
rect 255 -493 289 -459
rect 323 -493 357 -459
rect 391 -493 425 -459
rect 459 -493 493 -459
rect 527 -493 561 -459
rect 595 -493 629 -459
rect 663 -493 697 -459
rect 731 -493 765 -459
rect 799 -493 833 -459
rect 867 -493 901 -459
rect 935 -493 969 -459
rect 1003 -493 1037 -459
<< poly >>
rect -995 391 -925 407
rect -995 357 -977 391
rect -943 357 -925 391
rect -995 319 -925 357
rect -867 391 -797 407
rect -867 357 -849 391
rect -815 357 -797 391
rect -867 319 -797 357
rect -739 391 -669 407
rect -739 357 -721 391
rect -687 357 -669 391
rect -739 319 -669 357
rect -611 391 -541 407
rect -611 357 -593 391
rect -559 357 -541 391
rect -611 319 -541 357
rect -483 391 -413 407
rect -483 357 -465 391
rect -431 357 -413 391
rect -483 319 -413 357
rect -355 391 -285 407
rect -355 357 -337 391
rect -303 357 -285 391
rect -355 319 -285 357
rect -227 391 -157 407
rect -227 357 -209 391
rect -175 357 -157 391
rect -227 319 -157 357
rect -99 391 -29 407
rect -99 357 -81 391
rect -47 357 -29 391
rect -99 319 -29 357
rect 29 391 99 407
rect 29 357 47 391
rect 81 357 99 391
rect 29 319 99 357
rect 157 391 227 407
rect 157 357 175 391
rect 209 357 227 391
rect 157 319 227 357
rect 285 391 355 407
rect 285 357 303 391
rect 337 357 355 391
rect 285 319 355 357
rect 413 391 483 407
rect 413 357 431 391
rect 465 357 483 391
rect 413 319 483 357
rect 541 391 611 407
rect 541 357 559 391
rect 593 357 611 391
rect 541 319 611 357
rect 669 391 739 407
rect 669 357 687 391
rect 721 357 739 391
rect 669 319 739 357
rect 797 391 867 407
rect 797 357 815 391
rect 849 357 867 391
rect 797 319 867 357
rect 925 391 995 407
rect 925 357 943 391
rect 977 357 995 391
rect 925 319 995 357
rect -995 -407 -925 -381
rect -867 -407 -797 -381
rect -739 -407 -669 -381
rect -611 -407 -541 -381
rect -483 -407 -413 -381
rect -355 -407 -285 -381
rect -227 -407 -157 -381
rect -99 -407 -29 -381
rect 29 -407 99 -381
rect 157 -407 227 -381
rect 285 -407 355 -381
rect 413 -407 483 -381
rect 541 -407 611 -381
rect 669 -407 739 -381
rect 797 -407 867 -381
rect 925 -407 995 -381
<< polycont >>
rect -977 357 -943 391
rect -849 357 -815 391
rect -721 357 -687 391
rect -593 357 -559 391
rect -465 357 -431 391
rect -337 357 -303 391
rect -209 357 -175 391
rect -81 357 -47 391
rect 47 357 81 391
rect 175 357 209 391
rect 303 357 337 391
rect 431 357 465 391
rect 559 357 593 391
rect 687 357 721 391
rect 815 357 849 391
rect 943 357 977 391
<< locali >>
rect -1155 459 -1037 493
rect -1003 459 -969 493
rect -935 459 -901 493
rect -867 459 -833 493
rect -799 459 -765 493
rect -731 459 -697 493
rect -663 459 -629 493
rect -595 459 -561 493
rect -527 459 -493 493
rect -459 459 -425 493
rect -391 459 -357 493
rect -323 459 -289 493
rect -255 459 -221 493
rect -187 459 -153 493
rect -119 459 -85 493
rect -51 459 -17 493
rect 17 459 51 493
rect 85 459 119 493
rect 153 459 187 493
rect 221 459 255 493
rect 289 459 323 493
rect 357 459 391 493
rect 425 459 459 493
rect 493 459 527 493
rect 561 459 595 493
rect 629 459 663 493
rect 697 459 731 493
rect 765 459 799 493
rect 833 459 867 493
rect 901 459 935 493
rect 969 459 1003 493
rect 1037 459 1155 493
rect -1155 391 -1121 459
rect 1121 391 1155 459
rect -995 357 -977 391
rect -943 357 -925 391
rect -867 357 -849 391
rect -815 357 -797 391
rect -739 357 -721 391
rect -687 357 -669 391
rect -611 357 -593 391
rect -559 357 -541 391
rect -483 357 -465 391
rect -431 357 -413 391
rect -355 357 -337 391
rect -303 357 -285 391
rect -227 357 -209 391
rect -175 357 -157 391
rect -99 357 -81 391
rect -47 357 -29 391
rect 29 357 47 391
rect 81 357 99 391
rect 157 357 175 391
rect 209 357 227 391
rect 285 357 303 391
rect 337 357 355 391
rect 413 357 431 391
rect 465 357 483 391
rect 541 357 559 391
rect 593 357 611 391
rect 669 357 687 391
rect 721 357 739 391
rect 797 357 815 391
rect 849 357 867 391
rect 925 357 943 391
rect 977 357 995 391
rect -1155 323 -1121 357
rect 1121 323 1155 357
rect -1155 255 -1121 289
rect -1155 187 -1121 221
rect -1155 119 -1121 153
rect -1155 51 -1121 85
rect -1155 -17 -1121 17
rect -1155 -85 -1121 -51
rect -1155 -153 -1121 -119
rect -1155 -221 -1121 -187
rect -1155 -289 -1121 -255
rect -1155 -357 -1121 -323
rect -1041 292 -1007 323
rect -1041 224 -1007 240
rect -1041 156 -1007 168
rect -1041 88 -1007 96
rect -1041 20 -1007 24
rect -1041 -86 -1007 -82
rect -1041 -158 -1007 -150
rect -1041 -230 -1007 -218
rect -1041 -302 -1007 -286
rect -1041 -385 -1007 -354
rect -913 292 -879 323
rect -913 224 -879 240
rect -913 156 -879 168
rect -913 88 -879 96
rect -913 20 -879 24
rect -913 -86 -879 -82
rect -913 -158 -879 -150
rect -913 -230 -879 -218
rect -913 -302 -879 -286
rect -913 -385 -879 -354
rect -785 292 -751 323
rect -785 224 -751 240
rect -785 156 -751 168
rect -785 88 -751 96
rect -785 20 -751 24
rect -785 -86 -751 -82
rect -785 -158 -751 -150
rect -785 -230 -751 -218
rect -785 -302 -751 -286
rect -785 -385 -751 -354
rect -657 292 -623 323
rect -657 224 -623 240
rect -657 156 -623 168
rect -657 88 -623 96
rect -657 20 -623 24
rect -657 -86 -623 -82
rect -657 -158 -623 -150
rect -657 -230 -623 -218
rect -657 -302 -623 -286
rect -657 -385 -623 -354
rect -529 292 -495 323
rect -529 224 -495 240
rect -529 156 -495 168
rect -529 88 -495 96
rect -529 20 -495 24
rect -529 -86 -495 -82
rect -529 -158 -495 -150
rect -529 -230 -495 -218
rect -529 -302 -495 -286
rect -529 -385 -495 -354
rect -401 292 -367 323
rect -401 224 -367 240
rect -401 156 -367 168
rect -401 88 -367 96
rect -401 20 -367 24
rect -401 -86 -367 -82
rect -401 -158 -367 -150
rect -401 -230 -367 -218
rect -401 -302 -367 -286
rect -401 -385 -367 -354
rect -273 292 -239 323
rect -273 224 -239 240
rect -273 156 -239 168
rect -273 88 -239 96
rect -273 20 -239 24
rect -273 -86 -239 -82
rect -273 -158 -239 -150
rect -273 -230 -239 -218
rect -273 -302 -239 -286
rect -273 -385 -239 -354
rect -145 292 -111 323
rect -145 224 -111 240
rect -145 156 -111 168
rect -145 88 -111 96
rect -145 20 -111 24
rect -145 -86 -111 -82
rect -145 -158 -111 -150
rect -145 -230 -111 -218
rect -145 -302 -111 -286
rect -145 -385 -111 -354
rect -17 292 17 323
rect -17 224 17 240
rect -17 156 17 168
rect -17 88 17 96
rect -17 20 17 24
rect -17 -86 17 -82
rect -17 -158 17 -150
rect -17 -230 17 -218
rect -17 -302 17 -286
rect -17 -385 17 -354
rect 111 292 145 323
rect 111 224 145 240
rect 111 156 145 168
rect 111 88 145 96
rect 111 20 145 24
rect 111 -86 145 -82
rect 111 -158 145 -150
rect 111 -230 145 -218
rect 111 -302 145 -286
rect 111 -385 145 -354
rect 239 292 273 323
rect 239 224 273 240
rect 239 156 273 168
rect 239 88 273 96
rect 239 20 273 24
rect 239 -86 273 -82
rect 239 -158 273 -150
rect 239 -230 273 -218
rect 239 -302 273 -286
rect 239 -385 273 -354
rect 367 292 401 323
rect 367 224 401 240
rect 367 156 401 168
rect 367 88 401 96
rect 367 20 401 24
rect 367 -86 401 -82
rect 367 -158 401 -150
rect 367 -230 401 -218
rect 367 -302 401 -286
rect 367 -385 401 -354
rect 495 292 529 323
rect 495 224 529 240
rect 495 156 529 168
rect 495 88 529 96
rect 495 20 529 24
rect 495 -86 529 -82
rect 495 -158 529 -150
rect 495 -230 529 -218
rect 495 -302 529 -286
rect 495 -385 529 -354
rect 623 292 657 323
rect 623 224 657 240
rect 623 156 657 168
rect 623 88 657 96
rect 623 20 657 24
rect 623 -86 657 -82
rect 623 -158 657 -150
rect 623 -230 657 -218
rect 623 -302 657 -286
rect 623 -385 657 -354
rect 751 292 785 323
rect 751 224 785 240
rect 751 156 785 168
rect 751 88 785 96
rect 751 20 785 24
rect 751 -86 785 -82
rect 751 -158 785 -150
rect 751 -230 785 -218
rect 751 -302 785 -286
rect 751 -385 785 -354
rect 879 292 913 323
rect 879 224 913 240
rect 879 156 913 168
rect 879 88 913 96
rect 879 20 913 24
rect 879 -86 913 -82
rect 879 -158 913 -150
rect 879 -230 913 -218
rect 879 -302 913 -286
rect 879 -385 913 -354
rect 1007 292 1041 323
rect 1007 224 1041 240
rect 1007 156 1041 168
rect 1007 88 1041 96
rect 1007 20 1041 24
rect 1007 -86 1041 -82
rect 1007 -158 1041 -150
rect 1007 -230 1041 -218
rect 1007 -302 1041 -286
rect 1007 -385 1041 -354
rect 1121 255 1155 289
rect 1121 187 1155 221
rect 1121 119 1155 153
rect 1121 51 1155 85
rect 1121 -17 1155 17
rect 1121 -85 1155 -51
rect 1121 -153 1155 -119
rect 1121 -221 1155 -187
rect 1121 -289 1155 -255
rect 1121 -357 1155 -323
rect -1155 -459 -1121 -391
rect 1121 -459 1155 -391
rect -1155 -493 -1037 -459
rect -1003 -493 -969 -459
rect -935 -493 -901 -459
rect -867 -493 -833 -459
rect -799 -493 -765 -459
rect -731 -493 -697 -459
rect -663 -493 -629 -459
rect -595 -493 -561 -459
rect -527 -493 -493 -459
rect -459 -493 -425 -459
rect -391 -493 -357 -459
rect -323 -493 -289 -459
rect -255 -493 -221 -459
rect -187 -493 -153 -459
rect -119 -493 -85 -459
rect -51 -493 -17 -459
rect 17 -493 51 -459
rect 85 -493 119 -459
rect 153 -493 187 -459
rect 221 -493 255 -459
rect 289 -493 323 -459
rect 357 -493 391 -459
rect 425 -493 459 -459
rect 493 -493 527 -459
rect 561 -493 595 -459
rect 629 -493 663 -459
rect 697 -493 731 -459
rect 765 -493 799 -459
rect 833 -493 867 -459
rect 901 -493 935 -459
rect 969 -493 1003 -459
rect 1037 -493 1155 -459
<< viali >>
rect -977 357 -943 391
rect -849 357 -815 391
rect -721 357 -687 391
rect -593 357 -559 391
rect -465 357 -431 391
rect -337 357 -303 391
rect -209 357 -175 391
rect -81 357 -47 391
rect 47 357 81 391
rect 175 357 209 391
rect 303 357 337 391
rect 431 357 465 391
rect 559 357 593 391
rect 687 357 721 391
rect 815 357 849 391
rect 943 357 977 391
rect -1041 258 -1007 274
rect -1041 240 -1007 258
rect -1041 190 -1007 202
rect -1041 168 -1007 190
rect -1041 122 -1007 130
rect -1041 96 -1007 122
rect -1041 54 -1007 58
rect -1041 24 -1007 54
rect -1041 -48 -1007 -14
rect -1041 -116 -1007 -86
rect -1041 -120 -1007 -116
rect -1041 -184 -1007 -158
rect -1041 -192 -1007 -184
rect -1041 -252 -1007 -230
rect -1041 -264 -1007 -252
rect -1041 -320 -1007 -302
rect -1041 -336 -1007 -320
rect -913 258 -879 274
rect -913 240 -879 258
rect -913 190 -879 202
rect -913 168 -879 190
rect -913 122 -879 130
rect -913 96 -879 122
rect -913 54 -879 58
rect -913 24 -879 54
rect -913 -48 -879 -14
rect -913 -116 -879 -86
rect -913 -120 -879 -116
rect -913 -184 -879 -158
rect -913 -192 -879 -184
rect -913 -252 -879 -230
rect -913 -264 -879 -252
rect -913 -320 -879 -302
rect -913 -336 -879 -320
rect -785 258 -751 274
rect -785 240 -751 258
rect -785 190 -751 202
rect -785 168 -751 190
rect -785 122 -751 130
rect -785 96 -751 122
rect -785 54 -751 58
rect -785 24 -751 54
rect -785 -48 -751 -14
rect -785 -116 -751 -86
rect -785 -120 -751 -116
rect -785 -184 -751 -158
rect -785 -192 -751 -184
rect -785 -252 -751 -230
rect -785 -264 -751 -252
rect -785 -320 -751 -302
rect -785 -336 -751 -320
rect -657 258 -623 274
rect -657 240 -623 258
rect -657 190 -623 202
rect -657 168 -623 190
rect -657 122 -623 130
rect -657 96 -623 122
rect -657 54 -623 58
rect -657 24 -623 54
rect -657 -48 -623 -14
rect -657 -116 -623 -86
rect -657 -120 -623 -116
rect -657 -184 -623 -158
rect -657 -192 -623 -184
rect -657 -252 -623 -230
rect -657 -264 -623 -252
rect -657 -320 -623 -302
rect -657 -336 -623 -320
rect -529 258 -495 274
rect -529 240 -495 258
rect -529 190 -495 202
rect -529 168 -495 190
rect -529 122 -495 130
rect -529 96 -495 122
rect -529 54 -495 58
rect -529 24 -495 54
rect -529 -48 -495 -14
rect -529 -116 -495 -86
rect -529 -120 -495 -116
rect -529 -184 -495 -158
rect -529 -192 -495 -184
rect -529 -252 -495 -230
rect -529 -264 -495 -252
rect -529 -320 -495 -302
rect -529 -336 -495 -320
rect -401 258 -367 274
rect -401 240 -367 258
rect -401 190 -367 202
rect -401 168 -367 190
rect -401 122 -367 130
rect -401 96 -367 122
rect -401 54 -367 58
rect -401 24 -367 54
rect -401 -48 -367 -14
rect -401 -116 -367 -86
rect -401 -120 -367 -116
rect -401 -184 -367 -158
rect -401 -192 -367 -184
rect -401 -252 -367 -230
rect -401 -264 -367 -252
rect -401 -320 -367 -302
rect -401 -336 -367 -320
rect -273 258 -239 274
rect -273 240 -239 258
rect -273 190 -239 202
rect -273 168 -239 190
rect -273 122 -239 130
rect -273 96 -239 122
rect -273 54 -239 58
rect -273 24 -239 54
rect -273 -48 -239 -14
rect -273 -116 -239 -86
rect -273 -120 -239 -116
rect -273 -184 -239 -158
rect -273 -192 -239 -184
rect -273 -252 -239 -230
rect -273 -264 -239 -252
rect -273 -320 -239 -302
rect -273 -336 -239 -320
rect -145 258 -111 274
rect -145 240 -111 258
rect -145 190 -111 202
rect -145 168 -111 190
rect -145 122 -111 130
rect -145 96 -111 122
rect -145 54 -111 58
rect -145 24 -111 54
rect -145 -48 -111 -14
rect -145 -116 -111 -86
rect -145 -120 -111 -116
rect -145 -184 -111 -158
rect -145 -192 -111 -184
rect -145 -252 -111 -230
rect -145 -264 -111 -252
rect -145 -320 -111 -302
rect -145 -336 -111 -320
rect -17 258 17 274
rect -17 240 17 258
rect -17 190 17 202
rect -17 168 17 190
rect -17 122 17 130
rect -17 96 17 122
rect -17 54 17 58
rect -17 24 17 54
rect -17 -48 17 -14
rect -17 -116 17 -86
rect -17 -120 17 -116
rect -17 -184 17 -158
rect -17 -192 17 -184
rect -17 -252 17 -230
rect -17 -264 17 -252
rect -17 -320 17 -302
rect -17 -336 17 -320
rect 111 258 145 274
rect 111 240 145 258
rect 111 190 145 202
rect 111 168 145 190
rect 111 122 145 130
rect 111 96 145 122
rect 111 54 145 58
rect 111 24 145 54
rect 111 -48 145 -14
rect 111 -116 145 -86
rect 111 -120 145 -116
rect 111 -184 145 -158
rect 111 -192 145 -184
rect 111 -252 145 -230
rect 111 -264 145 -252
rect 111 -320 145 -302
rect 111 -336 145 -320
rect 239 258 273 274
rect 239 240 273 258
rect 239 190 273 202
rect 239 168 273 190
rect 239 122 273 130
rect 239 96 273 122
rect 239 54 273 58
rect 239 24 273 54
rect 239 -48 273 -14
rect 239 -116 273 -86
rect 239 -120 273 -116
rect 239 -184 273 -158
rect 239 -192 273 -184
rect 239 -252 273 -230
rect 239 -264 273 -252
rect 239 -320 273 -302
rect 239 -336 273 -320
rect 367 258 401 274
rect 367 240 401 258
rect 367 190 401 202
rect 367 168 401 190
rect 367 122 401 130
rect 367 96 401 122
rect 367 54 401 58
rect 367 24 401 54
rect 367 -48 401 -14
rect 367 -116 401 -86
rect 367 -120 401 -116
rect 367 -184 401 -158
rect 367 -192 401 -184
rect 367 -252 401 -230
rect 367 -264 401 -252
rect 367 -320 401 -302
rect 367 -336 401 -320
rect 495 258 529 274
rect 495 240 529 258
rect 495 190 529 202
rect 495 168 529 190
rect 495 122 529 130
rect 495 96 529 122
rect 495 54 529 58
rect 495 24 529 54
rect 495 -48 529 -14
rect 495 -116 529 -86
rect 495 -120 529 -116
rect 495 -184 529 -158
rect 495 -192 529 -184
rect 495 -252 529 -230
rect 495 -264 529 -252
rect 495 -320 529 -302
rect 495 -336 529 -320
rect 623 258 657 274
rect 623 240 657 258
rect 623 190 657 202
rect 623 168 657 190
rect 623 122 657 130
rect 623 96 657 122
rect 623 54 657 58
rect 623 24 657 54
rect 623 -48 657 -14
rect 623 -116 657 -86
rect 623 -120 657 -116
rect 623 -184 657 -158
rect 623 -192 657 -184
rect 623 -252 657 -230
rect 623 -264 657 -252
rect 623 -320 657 -302
rect 623 -336 657 -320
rect 751 258 785 274
rect 751 240 785 258
rect 751 190 785 202
rect 751 168 785 190
rect 751 122 785 130
rect 751 96 785 122
rect 751 54 785 58
rect 751 24 785 54
rect 751 -48 785 -14
rect 751 -116 785 -86
rect 751 -120 785 -116
rect 751 -184 785 -158
rect 751 -192 785 -184
rect 751 -252 785 -230
rect 751 -264 785 -252
rect 751 -320 785 -302
rect 751 -336 785 -320
rect 879 258 913 274
rect 879 240 913 258
rect 879 190 913 202
rect 879 168 913 190
rect 879 122 913 130
rect 879 96 913 122
rect 879 54 913 58
rect 879 24 913 54
rect 879 -48 913 -14
rect 879 -116 913 -86
rect 879 -120 913 -116
rect 879 -184 913 -158
rect 879 -192 913 -184
rect 879 -252 913 -230
rect 879 -264 913 -252
rect 879 -320 913 -302
rect 879 -336 913 -320
rect 1007 258 1041 274
rect 1007 240 1041 258
rect 1007 190 1041 202
rect 1007 168 1041 190
rect 1007 122 1041 130
rect 1007 96 1041 122
rect 1007 54 1041 58
rect 1007 24 1041 54
rect 1007 -48 1041 -14
rect 1007 -116 1041 -86
rect 1007 -120 1041 -116
rect 1007 -184 1041 -158
rect 1007 -192 1041 -184
rect 1007 -252 1041 -230
rect 1007 -264 1041 -252
rect 1007 -320 1041 -302
rect 1007 -336 1041 -320
<< metal1 >>
rect -991 391 -929 397
rect -991 357 -977 391
rect -943 357 -929 391
rect -991 351 -929 357
rect -863 391 -801 397
rect -863 357 -849 391
rect -815 357 -801 391
rect -863 351 -801 357
rect -735 391 -673 397
rect -735 357 -721 391
rect -687 357 -673 391
rect -735 351 -673 357
rect -607 391 -545 397
rect -607 357 -593 391
rect -559 357 -545 391
rect -607 351 -545 357
rect -479 391 -417 397
rect -479 357 -465 391
rect -431 357 -417 391
rect -479 351 -417 357
rect -351 391 -289 397
rect -351 357 -337 391
rect -303 357 -289 391
rect -351 351 -289 357
rect -223 391 -161 397
rect -223 357 -209 391
rect -175 357 -161 391
rect -223 351 -161 357
rect -95 391 -33 397
rect -95 357 -81 391
rect -47 357 -33 391
rect -95 351 -33 357
rect 33 391 95 397
rect 33 357 47 391
rect 81 357 95 391
rect 33 351 95 357
rect 161 391 223 397
rect 161 357 175 391
rect 209 357 223 391
rect 161 351 223 357
rect 289 391 351 397
rect 289 357 303 391
rect 337 357 351 391
rect 289 351 351 357
rect 417 391 479 397
rect 417 357 431 391
rect 465 357 479 391
rect 417 351 479 357
rect 545 391 607 397
rect 545 357 559 391
rect 593 357 607 391
rect 545 351 607 357
rect 673 391 735 397
rect 673 357 687 391
rect 721 357 735 391
rect 673 351 735 357
rect 801 391 863 397
rect 801 357 815 391
rect 849 357 863 391
rect 801 351 863 357
rect 929 391 991 397
rect 929 357 943 391
rect 977 357 991 391
rect 929 351 991 357
rect -1047 274 -1001 319
rect -1047 240 -1041 274
rect -1007 240 -1001 274
rect -1047 202 -1001 240
rect -1047 168 -1041 202
rect -1007 168 -1001 202
rect -1047 130 -1001 168
rect -1047 96 -1041 130
rect -1007 96 -1001 130
rect -1047 58 -1001 96
rect -1047 24 -1041 58
rect -1007 24 -1001 58
rect -1047 -14 -1001 24
rect -1047 -48 -1041 -14
rect -1007 -48 -1001 -14
rect -1047 -86 -1001 -48
rect -1047 -120 -1041 -86
rect -1007 -120 -1001 -86
rect -1047 -158 -1001 -120
rect -1047 -192 -1041 -158
rect -1007 -192 -1001 -158
rect -1047 -230 -1001 -192
rect -1047 -264 -1041 -230
rect -1007 -264 -1001 -230
rect -1047 -302 -1001 -264
rect -1047 -336 -1041 -302
rect -1007 -336 -1001 -302
rect -1047 -381 -1001 -336
rect -919 274 -873 319
rect -919 240 -913 274
rect -879 240 -873 274
rect -919 202 -873 240
rect -919 168 -913 202
rect -879 168 -873 202
rect -919 130 -873 168
rect -919 96 -913 130
rect -879 96 -873 130
rect -919 58 -873 96
rect -919 24 -913 58
rect -879 24 -873 58
rect -919 -14 -873 24
rect -919 -48 -913 -14
rect -879 -48 -873 -14
rect -919 -86 -873 -48
rect -919 -120 -913 -86
rect -879 -120 -873 -86
rect -919 -158 -873 -120
rect -919 -192 -913 -158
rect -879 -192 -873 -158
rect -919 -230 -873 -192
rect -919 -264 -913 -230
rect -879 -264 -873 -230
rect -919 -302 -873 -264
rect -919 -336 -913 -302
rect -879 -336 -873 -302
rect -919 -381 -873 -336
rect -791 274 -745 319
rect -791 240 -785 274
rect -751 240 -745 274
rect -791 202 -745 240
rect -791 168 -785 202
rect -751 168 -745 202
rect -791 130 -745 168
rect -791 96 -785 130
rect -751 96 -745 130
rect -791 58 -745 96
rect -791 24 -785 58
rect -751 24 -745 58
rect -791 -14 -745 24
rect -791 -48 -785 -14
rect -751 -48 -745 -14
rect -791 -86 -745 -48
rect -791 -120 -785 -86
rect -751 -120 -745 -86
rect -791 -158 -745 -120
rect -791 -192 -785 -158
rect -751 -192 -745 -158
rect -791 -230 -745 -192
rect -791 -264 -785 -230
rect -751 -264 -745 -230
rect -791 -302 -745 -264
rect -791 -336 -785 -302
rect -751 -336 -745 -302
rect -791 -381 -745 -336
rect -663 274 -617 319
rect -663 240 -657 274
rect -623 240 -617 274
rect -663 202 -617 240
rect -663 168 -657 202
rect -623 168 -617 202
rect -663 130 -617 168
rect -663 96 -657 130
rect -623 96 -617 130
rect -663 58 -617 96
rect -663 24 -657 58
rect -623 24 -617 58
rect -663 -14 -617 24
rect -663 -48 -657 -14
rect -623 -48 -617 -14
rect -663 -86 -617 -48
rect -663 -120 -657 -86
rect -623 -120 -617 -86
rect -663 -158 -617 -120
rect -663 -192 -657 -158
rect -623 -192 -617 -158
rect -663 -230 -617 -192
rect -663 -264 -657 -230
rect -623 -264 -617 -230
rect -663 -302 -617 -264
rect -663 -336 -657 -302
rect -623 -336 -617 -302
rect -663 -381 -617 -336
rect -535 274 -489 319
rect -535 240 -529 274
rect -495 240 -489 274
rect -535 202 -489 240
rect -535 168 -529 202
rect -495 168 -489 202
rect -535 130 -489 168
rect -535 96 -529 130
rect -495 96 -489 130
rect -535 58 -489 96
rect -535 24 -529 58
rect -495 24 -489 58
rect -535 -14 -489 24
rect -535 -48 -529 -14
rect -495 -48 -489 -14
rect -535 -86 -489 -48
rect -535 -120 -529 -86
rect -495 -120 -489 -86
rect -535 -158 -489 -120
rect -535 -192 -529 -158
rect -495 -192 -489 -158
rect -535 -230 -489 -192
rect -535 -264 -529 -230
rect -495 -264 -489 -230
rect -535 -302 -489 -264
rect -535 -336 -529 -302
rect -495 -336 -489 -302
rect -535 -381 -489 -336
rect -407 274 -361 319
rect -407 240 -401 274
rect -367 240 -361 274
rect -407 202 -361 240
rect -407 168 -401 202
rect -367 168 -361 202
rect -407 130 -361 168
rect -407 96 -401 130
rect -367 96 -361 130
rect -407 58 -361 96
rect -407 24 -401 58
rect -367 24 -361 58
rect -407 -14 -361 24
rect -407 -48 -401 -14
rect -367 -48 -361 -14
rect -407 -86 -361 -48
rect -407 -120 -401 -86
rect -367 -120 -361 -86
rect -407 -158 -361 -120
rect -407 -192 -401 -158
rect -367 -192 -361 -158
rect -407 -230 -361 -192
rect -407 -264 -401 -230
rect -367 -264 -361 -230
rect -407 -302 -361 -264
rect -407 -336 -401 -302
rect -367 -336 -361 -302
rect -407 -381 -361 -336
rect -279 274 -233 319
rect -279 240 -273 274
rect -239 240 -233 274
rect -279 202 -233 240
rect -279 168 -273 202
rect -239 168 -233 202
rect -279 130 -233 168
rect -279 96 -273 130
rect -239 96 -233 130
rect -279 58 -233 96
rect -279 24 -273 58
rect -239 24 -233 58
rect -279 -14 -233 24
rect -279 -48 -273 -14
rect -239 -48 -233 -14
rect -279 -86 -233 -48
rect -279 -120 -273 -86
rect -239 -120 -233 -86
rect -279 -158 -233 -120
rect -279 -192 -273 -158
rect -239 -192 -233 -158
rect -279 -230 -233 -192
rect -279 -264 -273 -230
rect -239 -264 -233 -230
rect -279 -302 -233 -264
rect -279 -336 -273 -302
rect -239 -336 -233 -302
rect -279 -381 -233 -336
rect -151 274 -105 319
rect -151 240 -145 274
rect -111 240 -105 274
rect -151 202 -105 240
rect -151 168 -145 202
rect -111 168 -105 202
rect -151 130 -105 168
rect -151 96 -145 130
rect -111 96 -105 130
rect -151 58 -105 96
rect -151 24 -145 58
rect -111 24 -105 58
rect -151 -14 -105 24
rect -151 -48 -145 -14
rect -111 -48 -105 -14
rect -151 -86 -105 -48
rect -151 -120 -145 -86
rect -111 -120 -105 -86
rect -151 -158 -105 -120
rect -151 -192 -145 -158
rect -111 -192 -105 -158
rect -151 -230 -105 -192
rect -151 -264 -145 -230
rect -111 -264 -105 -230
rect -151 -302 -105 -264
rect -151 -336 -145 -302
rect -111 -336 -105 -302
rect -151 -381 -105 -336
rect -23 274 23 319
rect -23 240 -17 274
rect 17 240 23 274
rect -23 202 23 240
rect -23 168 -17 202
rect 17 168 23 202
rect -23 130 23 168
rect -23 96 -17 130
rect 17 96 23 130
rect -23 58 23 96
rect -23 24 -17 58
rect 17 24 23 58
rect -23 -14 23 24
rect -23 -48 -17 -14
rect 17 -48 23 -14
rect -23 -86 23 -48
rect -23 -120 -17 -86
rect 17 -120 23 -86
rect -23 -158 23 -120
rect -23 -192 -17 -158
rect 17 -192 23 -158
rect -23 -230 23 -192
rect -23 -264 -17 -230
rect 17 -264 23 -230
rect -23 -302 23 -264
rect -23 -336 -17 -302
rect 17 -336 23 -302
rect -23 -381 23 -336
rect 105 274 151 319
rect 105 240 111 274
rect 145 240 151 274
rect 105 202 151 240
rect 105 168 111 202
rect 145 168 151 202
rect 105 130 151 168
rect 105 96 111 130
rect 145 96 151 130
rect 105 58 151 96
rect 105 24 111 58
rect 145 24 151 58
rect 105 -14 151 24
rect 105 -48 111 -14
rect 145 -48 151 -14
rect 105 -86 151 -48
rect 105 -120 111 -86
rect 145 -120 151 -86
rect 105 -158 151 -120
rect 105 -192 111 -158
rect 145 -192 151 -158
rect 105 -230 151 -192
rect 105 -264 111 -230
rect 145 -264 151 -230
rect 105 -302 151 -264
rect 105 -336 111 -302
rect 145 -336 151 -302
rect 105 -381 151 -336
rect 233 274 279 319
rect 233 240 239 274
rect 273 240 279 274
rect 233 202 279 240
rect 233 168 239 202
rect 273 168 279 202
rect 233 130 279 168
rect 233 96 239 130
rect 273 96 279 130
rect 233 58 279 96
rect 233 24 239 58
rect 273 24 279 58
rect 233 -14 279 24
rect 233 -48 239 -14
rect 273 -48 279 -14
rect 233 -86 279 -48
rect 233 -120 239 -86
rect 273 -120 279 -86
rect 233 -158 279 -120
rect 233 -192 239 -158
rect 273 -192 279 -158
rect 233 -230 279 -192
rect 233 -264 239 -230
rect 273 -264 279 -230
rect 233 -302 279 -264
rect 233 -336 239 -302
rect 273 -336 279 -302
rect 233 -381 279 -336
rect 361 274 407 319
rect 361 240 367 274
rect 401 240 407 274
rect 361 202 407 240
rect 361 168 367 202
rect 401 168 407 202
rect 361 130 407 168
rect 361 96 367 130
rect 401 96 407 130
rect 361 58 407 96
rect 361 24 367 58
rect 401 24 407 58
rect 361 -14 407 24
rect 361 -48 367 -14
rect 401 -48 407 -14
rect 361 -86 407 -48
rect 361 -120 367 -86
rect 401 -120 407 -86
rect 361 -158 407 -120
rect 361 -192 367 -158
rect 401 -192 407 -158
rect 361 -230 407 -192
rect 361 -264 367 -230
rect 401 -264 407 -230
rect 361 -302 407 -264
rect 361 -336 367 -302
rect 401 -336 407 -302
rect 361 -381 407 -336
rect 489 274 535 319
rect 489 240 495 274
rect 529 240 535 274
rect 489 202 535 240
rect 489 168 495 202
rect 529 168 535 202
rect 489 130 535 168
rect 489 96 495 130
rect 529 96 535 130
rect 489 58 535 96
rect 489 24 495 58
rect 529 24 535 58
rect 489 -14 535 24
rect 489 -48 495 -14
rect 529 -48 535 -14
rect 489 -86 535 -48
rect 489 -120 495 -86
rect 529 -120 535 -86
rect 489 -158 535 -120
rect 489 -192 495 -158
rect 529 -192 535 -158
rect 489 -230 535 -192
rect 489 -264 495 -230
rect 529 -264 535 -230
rect 489 -302 535 -264
rect 489 -336 495 -302
rect 529 -336 535 -302
rect 489 -381 535 -336
rect 617 274 663 319
rect 617 240 623 274
rect 657 240 663 274
rect 617 202 663 240
rect 617 168 623 202
rect 657 168 663 202
rect 617 130 663 168
rect 617 96 623 130
rect 657 96 663 130
rect 617 58 663 96
rect 617 24 623 58
rect 657 24 663 58
rect 617 -14 663 24
rect 617 -48 623 -14
rect 657 -48 663 -14
rect 617 -86 663 -48
rect 617 -120 623 -86
rect 657 -120 663 -86
rect 617 -158 663 -120
rect 617 -192 623 -158
rect 657 -192 663 -158
rect 617 -230 663 -192
rect 617 -264 623 -230
rect 657 -264 663 -230
rect 617 -302 663 -264
rect 617 -336 623 -302
rect 657 -336 663 -302
rect 617 -381 663 -336
rect 745 274 791 319
rect 745 240 751 274
rect 785 240 791 274
rect 745 202 791 240
rect 745 168 751 202
rect 785 168 791 202
rect 745 130 791 168
rect 745 96 751 130
rect 785 96 791 130
rect 745 58 791 96
rect 745 24 751 58
rect 785 24 791 58
rect 745 -14 791 24
rect 745 -48 751 -14
rect 785 -48 791 -14
rect 745 -86 791 -48
rect 745 -120 751 -86
rect 785 -120 791 -86
rect 745 -158 791 -120
rect 745 -192 751 -158
rect 785 -192 791 -158
rect 745 -230 791 -192
rect 745 -264 751 -230
rect 785 -264 791 -230
rect 745 -302 791 -264
rect 745 -336 751 -302
rect 785 -336 791 -302
rect 745 -381 791 -336
rect 873 274 919 319
rect 873 240 879 274
rect 913 240 919 274
rect 873 202 919 240
rect 873 168 879 202
rect 913 168 919 202
rect 873 130 919 168
rect 873 96 879 130
rect 913 96 919 130
rect 873 58 919 96
rect 873 24 879 58
rect 913 24 919 58
rect 873 -14 919 24
rect 873 -48 879 -14
rect 913 -48 919 -14
rect 873 -86 919 -48
rect 873 -120 879 -86
rect 913 -120 919 -86
rect 873 -158 919 -120
rect 873 -192 879 -158
rect 913 -192 919 -158
rect 873 -230 919 -192
rect 873 -264 879 -230
rect 913 -264 919 -230
rect 873 -302 919 -264
rect 873 -336 879 -302
rect 913 -336 919 -302
rect 873 -381 919 -336
rect 1001 274 1047 319
rect 1001 240 1007 274
rect 1041 240 1047 274
rect 1001 202 1047 240
rect 1001 168 1007 202
rect 1041 168 1047 202
rect 1001 130 1047 168
rect 1001 96 1007 130
rect 1041 96 1047 130
rect 1001 58 1047 96
rect 1001 24 1007 58
rect 1041 24 1047 58
rect 1001 -14 1047 24
rect 1001 -48 1007 -14
rect 1041 -48 1047 -14
rect 1001 -86 1047 -48
rect 1001 -120 1007 -86
rect 1041 -120 1047 -86
rect 1001 -158 1047 -120
rect 1001 -192 1007 -158
rect 1041 -192 1047 -158
rect 1001 -230 1047 -192
rect 1001 -264 1007 -230
rect 1041 -264 1047 -230
rect 1001 -302 1047 -264
rect 1001 -336 1007 -302
rect 1041 -336 1047 -302
rect 1001 -381 1047 -336
<< labels >>
flabel metal1 s -960 374 -960 374 0 FreeSans 300 0 0 0 G
port 1 nsew
flabel metal1 s -832 374 -832 374 0 FreeSans 300 0 0 0 G
port 1 nsew
flabel metal1 s -704 374 -704 374 0 FreeSans 300 0 0 0 G
port 1 nsew
flabel metal1 s -576 374 -576 374 0 FreeSans 300 0 0 0 G
port 1 nsew
flabel metal1 s -448 374 -448 374 0 FreeSans 300 0 0 0 G
port 1 nsew
flabel metal1 s -320 374 -320 374 0 FreeSans 300 0 0 0 G
port 1 nsew
flabel metal1 s -192 374 -192 374 0 FreeSans 300 0 0 0 G
port 1 nsew
flabel metal1 s -64 374 -64 374 0 FreeSans 300 0 0 0 G
port 1 nsew
flabel metal1 s 64 374 64 374 0 FreeSans 300 0 0 0 G
port 1 nsew
flabel metal1 s 192 374 192 374 0 FreeSans 300 0 0 0 G
port 1 nsew
flabel metal1 s 320 374 320 374 0 FreeSans 300 0 0 0 G
port 1 nsew
flabel metal1 s 448 374 448 374 0 FreeSans 300 0 0 0 G
port 1 nsew
flabel metal1 s 576 374 576 374 0 FreeSans 300 0 0 0 G
port 1 nsew
flabel metal1 s 704 374 704 374 0 FreeSans 300 0 0 0 G
port 1 nsew
flabel metal1 s 832 374 832 374 0 FreeSans 300 0 0 0 G
port 1 nsew
flabel metal1 s 960 374 960 374 0 FreeSans 300 0 0 0 G
port 1 nsew
flabel metal1 s -1024 -31 -1024 -31 0 FreeSans 300 0 0 0 D
port 2 nsew
flabel metal1 s -896 -31 -896 -31 0 FreeSans 300 0 0 0 S
port 3 nsew
flabel metal1 s -768 -31 -768 -31 0 FreeSans 300 0 0 0 D
port 2 nsew
flabel metal1 s -640 -31 -640 -31 0 FreeSans 300 0 0 0 S
port 3 nsew
flabel metal1 s -512 -31 -512 -31 0 FreeSans 300 0 0 0 D
port 2 nsew
flabel metal1 s -384 -31 -384 -31 0 FreeSans 300 0 0 0 S
port 3 nsew
flabel metal1 s -256 -31 -256 -31 0 FreeSans 300 0 0 0 D
port 2 nsew
flabel metal1 s -128 -31 -128 -31 0 FreeSans 300 0 0 0 S
port 3 nsew
flabel metal1 s 0 -31 0 -31 0 FreeSans 300 0 0 0 D
port 2 nsew
flabel metal1 s 128 -31 128 -31 0 FreeSans 300 0 0 0 S
port 3 nsew
flabel metal1 s 256 -31 256 -31 0 FreeSans 300 0 0 0 D
port 2 nsew
flabel metal1 s 384 -31 384 -31 0 FreeSans 300 0 0 0 S
port 3 nsew
flabel metal1 s 512 -31 512 -31 0 FreeSans 300 0 0 0 D
port 2 nsew
flabel metal1 s 640 -31 640 -31 0 FreeSans 300 0 0 0 S
port 3 nsew
flabel metal1 s 768 -31 768 -31 0 FreeSans 300 0 0 0 D
port 2 nsew
flabel metal1 s 896 -31 896 -31 0 FreeSans 300 0 0 0 S
port 3 nsew
flabel metal1 s 1024 -31 1024 -31 0 FreeSans 300 0 0 0 D
port 2 nsew
<< properties >>
string FIXED_BBOX -1138 -476 1138 476
<< end >>
