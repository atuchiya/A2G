magic
tech sky130A
magscale 1 2
timestamp 1680003372
<< viali >>
rect 1344 2878 1378 2912
rect 3620 2878 3654 2912
rect 4120 2878 4154 2912
rect 8444 2878 8478 2912
rect 8944 2878 8978 2912
rect 11220 2878 11254 2912
rect 1344 2806 1378 2840
rect 3620 2806 3654 2840
rect 4120 2806 4154 2840
rect 8444 2806 8478 2840
rect 8944 2806 8978 2840
rect 11220 2806 11254 2840
rect 1344 2734 1378 2768
rect 3620 2734 3654 2768
rect 4120 2734 4154 2768
rect 8444 2734 8478 2768
rect 8944 2734 8978 2768
rect 11220 2734 11254 2768
rect 1344 2662 1378 2696
rect 3620 2662 3654 2696
rect 4120 2662 4154 2696
rect 8444 2662 8478 2696
rect 8944 2662 8978 2696
rect 11220 2662 11254 2696
rect 1344 2590 1378 2624
rect 3620 2590 3654 2624
rect 4120 2590 4154 2624
rect 8444 2590 8478 2624
rect 8944 2590 8978 2624
rect 11220 2590 11254 2624
rect 1344 2518 1378 2552
rect 3620 2518 3654 2552
rect 4120 2518 4154 2552
rect 8444 2518 8478 2552
rect 8944 2518 8978 2552
rect 11220 2518 11254 2552
rect 1344 2446 1378 2480
rect 3620 2446 3654 2480
rect 4120 2446 4154 2480
rect 8444 2446 8478 2480
rect 8944 2446 8978 2480
rect 11220 2446 11254 2480
rect 1344 2374 1378 2408
rect 3620 2374 3654 2408
rect 4120 2374 4154 2408
rect 8444 2374 8478 2408
rect 8944 2374 8978 2408
rect 11220 2374 11254 2408
rect 1344 2302 1378 2336
rect 3620 2302 3654 2336
rect 4120 2302 4154 2336
rect 8444 2302 8478 2336
rect 8944 2302 8978 2336
rect 11220 2302 11254 2336
rect 1344 2230 1378 2264
rect 3620 2230 3654 2264
rect 4120 2230 4154 2264
rect 8444 2230 8478 2264
rect 8944 2230 8978 2264
rect 11220 2230 11254 2264
rect 1344 2158 1378 2192
rect 3620 2158 3654 2192
rect 4120 2158 4154 2192
rect 8444 2158 8478 2192
rect 8944 2158 8978 2192
rect 11220 2158 11254 2192
rect 1344 2086 1378 2120
rect 3620 2086 3654 2120
rect 4120 2086 4154 2120
rect 8444 2086 8478 2120
rect 8944 2086 8978 2120
rect 11220 2086 11254 2120
rect 408 1278 442 1312
rect 5756 1278 5790 1312
rect 6608 1278 6642 1312
rect 11956 1278 11990 1312
rect 408 1206 442 1240
rect 5756 1206 5790 1240
rect 6608 1206 6642 1240
rect 11956 1206 11990 1240
rect 408 1134 442 1168
rect 5756 1134 5790 1168
rect 6608 1134 6642 1168
rect 11956 1134 11990 1168
rect 408 1062 442 1096
rect 5756 1062 5790 1096
rect 6608 1062 6642 1096
rect 11956 1062 11990 1096
rect 408 990 442 1024
rect 5756 990 5790 1024
rect 6608 990 6642 1024
rect 11956 990 11990 1024
rect 408 918 442 952
rect 5756 918 5790 952
rect 6608 918 6642 952
rect 11956 918 11990 952
rect 408 846 442 880
rect 5756 846 5790 880
rect 6608 846 6642 880
rect 11956 846 11990 880
rect 408 774 442 808
rect 5756 774 5790 808
rect 6608 774 6642 808
rect 11956 774 11990 808
rect 408 702 442 736
rect 5756 702 5790 736
rect 6608 702 6642 736
rect 11956 702 11990 736
rect 408 630 442 664
rect 5756 630 5790 664
rect 6608 630 6642 664
rect 11956 630 11990 664
rect 408 558 442 592
rect 5756 558 5790 592
rect 6608 558 6642 592
rect 11956 558 11990 592
rect 408 486 442 520
rect 5756 486 5790 520
rect 6608 486 6642 520
rect 11956 486 11990 520
<< metal1 >>
rect -150 3550 -50 3600
rect 50 3550 150 3600
rect 250 3550 350 3600
rect 450 3550 550 3600
rect 650 3550 750 3600
rect 850 3550 950 3600
rect 1050 3550 1150 3600
rect 1250 3550 1350 3600
rect 1450 3550 1550 3600
rect 1650 3550 1750 3600
rect 1850 3550 1950 3600
rect 2050 3550 2150 3600
rect 2250 3550 2350 3600
rect 2450 3550 2550 3600
rect 2650 3550 2750 3600
rect 2850 3550 2950 3600
rect 3050 3550 3150 3600
rect 3250 3550 3350 3600
rect 3450 3550 3550 3600
rect 3650 3550 3750 3600
rect 3850 3550 3950 3600
rect 4050 3550 4150 3600
rect 4250 3550 4350 3600
rect 4450 3550 4550 3600
rect 4650 3550 4750 3600
rect 4850 3550 4950 3600
rect 5050 3550 5150 3600
rect 5250 3550 5350 3600
rect 5450 3550 5550 3600
rect 5650 3550 5750 3600
rect 5850 3550 5950 3600
rect 6050 3550 6150 3600
rect 6250 3550 6350 3600
rect 6450 3550 6550 3600
rect 6650 3550 6750 3600
rect 6850 3550 6950 3600
rect 7050 3550 7150 3600
rect 7250 3550 7350 3600
rect 7450 3550 7550 3600
rect 7650 3550 7750 3600
rect 7850 3550 7950 3600
rect 8050 3550 8150 3600
rect 8250 3550 8350 3600
rect 8450 3550 8550 3600
rect 8650 3550 8750 3600
rect 8850 3550 8950 3600
rect 9050 3550 9150 3600
rect 9250 3550 9350 3600
rect 9450 3550 9550 3600
rect 9650 3550 9750 3600
rect 9850 3550 9950 3600
rect 10050 3550 10150 3600
rect 10250 3550 10350 3600
rect 10450 3550 10550 3600
rect 10650 3550 10750 3600
rect 10850 3550 10950 3600
rect 11050 3550 11150 3600
rect 11250 3550 11350 3600
rect 11450 3550 11550 3600
rect 11650 3550 11750 3600
rect 11850 3550 11950 3600
rect 12050 3550 12150 3600
rect 12250 3550 12350 3600
rect 12450 3550 12550 3600
rect -200 3450 12600 3550
rect -150 3350 -50 3450
rect 50 3350 150 3450
rect 250 3350 350 3450
rect 450 3350 550 3450
rect 650 3350 750 3450
rect 850 3350 950 3450
rect 1050 3350 1150 3450
rect 1250 3350 1350 3450
rect 1450 3350 1550 3450
rect 1650 3350 1750 3450
rect 1850 3350 1950 3450
rect 2050 3350 2150 3450
rect 2250 3350 2350 3450
rect 2450 3350 2550 3450
rect 2650 3350 2750 3450
rect 2850 3350 2950 3450
rect 3050 3350 3150 3450
rect 3250 3350 3350 3450
rect 3450 3350 3550 3450
rect 3650 3350 3750 3450
rect 3850 3350 3950 3450
rect 4050 3350 4150 3450
rect 4250 3350 4350 3450
rect 4450 3350 4550 3450
rect 4650 3350 4750 3450
rect 4850 3350 4950 3450
rect 5050 3350 5150 3450
rect 5250 3350 5350 3450
rect 5450 3350 5550 3450
rect 5650 3350 5750 3450
rect 5850 3350 5950 3450
rect 6050 3350 6150 3450
rect 6250 3350 6350 3450
rect 6450 3350 6550 3450
rect 6650 3350 6750 3450
rect 6850 3350 6950 3450
rect 7050 3350 7150 3450
rect 7250 3350 7350 3450
rect 7450 3350 7550 3450
rect 7650 3350 7750 3450
rect 7850 3350 7950 3450
rect 8050 3350 8150 3450
rect 8250 3350 8350 3450
rect 8450 3350 8550 3450
rect 8650 3350 8750 3450
rect 8850 3350 8950 3450
rect 9050 3350 9150 3450
rect 9250 3350 9350 3450
rect 9450 3350 9550 3450
rect 9650 3350 9750 3450
rect 9850 3350 9950 3450
rect 10050 3350 10150 3450
rect 10250 3350 10350 3450
rect 10450 3350 10550 3450
rect 10650 3350 10750 3450
rect 10850 3350 10950 3450
rect 11050 3350 11150 3450
rect 11250 3350 11350 3450
rect 11450 3350 11550 3450
rect 11650 3350 11750 3450
rect 11850 3350 11950 3450
rect 12050 3350 12150 3450
rect 12250 3350 12350 3450
rect 12450 3350 12550 3450
rect -200 3250 12600 3350
rect -150 3150 -50 3250
rect 50 3150 150 3250
rect 250 3150 350 3250
rect 450 3150 550 3250
rect 650 3150 750 3250
rect 850 3150 950 3250
rect 1050 3150 1150 3250
rect 1250 3200 1350 3250
rect 1450 3200 1550 3250
rect 1650 3200 1750 3250
rect 1850 3200 1950 3250
rect 2050 3200 2150 3250
rect 2250 3200 2350 3250
rect 2450 3200 2550 3250
rect 2650 3200 2750 3250
rect 2850 3200 2950 3250
rect 3050 3200 3150 3250
rect 3250 3200 3350 3250
rect 3450 3200 3550 3250
rect 3650 3200 3750 3250
rect 3850 3150 3950 3250
rect 4050 3200 4150 3250
rect 4250 3200 4350 3250
rect 4450 3200 4550 3250
rect 4650 3200 4750 3250
rect 4850 3200 4950 3250
rect 5050 3200 5150 3250
rect 5250 3200 5350 3250
rect 5450 3200 5550 3250
rect 5650 3200 5750 3250
rect 5850 3200 5950 3250
rect 6050 3200 6150 3250
rect 6250 3200 6350 3250
rect 6450 3200 6550 3250
rect 6650 3200 6750 3250
rect 6850 3200 6950 3250
rect 7050 3200 7150 3250
rect 7250 3200 7350 3250
rect 7450 3200 7550 3250
rect 7650 3200 7750 3250
rect 7850 3200 7950 3250
rect 8050 3200 8150 3250
rect 8250 3200 8350 3250
rect 8450 3200 8550 3250
rect 8650 3150 8750 3250
rect 8850 3200 8950 3250
rect 9050 3200 9150 3250
rect 9250 3200 9350 3250
rect 9450 3200 9550 3250
rect 9650 3200 9750 3250
rect 9850 3200 9950 3250
rect 10050 3200 10150 3250
rect 10250 3200 10350 3250
rect 10450 3200 10550 3250
rect 10650 3200 10750 3250
rect 10850 3200 10950 3250
rect 11050 3200 11150 3250
rect 11250 3200 11350 3250
rect 11450 3150 11550 3250
rect 11650 3150 11750 3250
rect 11850 3150 11950 3250
rect 12050 3150 12150 3250
rect 12250 3150 12350 3250
rect 12450 3150 12550 3250
rect -200 3050 1200 3150
rect 3800 3050 4000 3150
rect 8600 3050 8800 3150
rect 11400 3050 12600 3150
rect -150 2950 -50 3050
rect 50 2950 150 3050
rect 250 2950 350 3050
rect 450 2950 550 3050
rect 650 2950 750 3050
rect 850 2950 950 3050
rect 1050 2950 1150 3050
rect -200 2850 1200 2950
rect 1322 2912 1402 2958
rect 1322 2878 1344 2912
rect 1378 2878 1402 2912
rect -150 2750 -50 2850
rect 50 2750 150 2850
rect 250 2750 350 2850
rect 450 2750 550 2850
rect 650 2750 750 2850
rect 850 2750 950 2850
rect 1050 2750 1150 2850
rect 1322 2840 1402 2878
rect 1322 2806 1344 2840
rect 1378 2806 1402 2840
rect 1322 2768 1402 2806
rect -200 2650 1200 2750
rect 1322 2734 1344 2768
rect 1378 2734 1402 2768
rect 1322 2696 1402 2734
rect 1322 2662 1344 2696
rect 1378 2662 1402 2696
rect -150 2550 -50 2650
rect 50 2550 150 2650
rect 250 2550 350 2650
rect 450 2550 550 2650
rect 650 2550 750 2650
rect 850 2550 950 2650
rect 1050 2550 1150 2650
rect 1322 2624 1402 2662
rect 1322 2590 1344 2624
rect 1378 2590 1402 2624
rect 1322 2552 1402 2590
rect -200 2450 1200 2550
rect 1322 2518 1344 2552
rect 1378 2518 1402 2552
rect 1322 2480 1402 2518
rect -150 2350 -50 2450
rect 50 2350 150 2450
rect 250 2350 350 2450
rect 450 2350 550 2450
rect 650 2350 750 2450
rect 850 2350 950 2450
rect 1050 2350 1150 2450
rect 1322 2446 1344 2480
rect 1378 2446 1402 2480
rect 1322 2408 1402 2446
rect 1322 2374 1344 2408
rect 1378 2374 1402 2408
rect -200 2250 1200 2350
rect 1322 2336 1402 2374
rect 1322 2302 1344 2336
rect 1378 2302 1402 2336
rect 1322 2264 1402 2302
rect -150 2150 -50 2250
rect 50 2150 150 2250
rect 250 2150 350 2250
rect 450 2150 550 2250
rect 650 2150 750 2250
rect 850 2150 950 2250
rect 1050 2150 1150 2250
rect 1322 2230 1344 2264
rect 1378 2230 1402 2264
rect 1322 2192 1402 2230
rect 1322 2158 1344 2192
rect 1378 2158 1402 2192
rect -200 2050 1200 2150
rect 1322 2120 1402 2158
rect 1322 2086 1344 2120
rect 1378 2086 1402 2120
rect -150 1950 -50 2050
rect 50 1950 150 2050
rect 250 1950 350 2050
rect 450 1950 550 2050
rect 650 1950 750 2050
rect 850 1950 950 2050
rect 1050 1950 1150 2050
rect 1322 2040 1402 2086
rect 3598 2912 3678 2958
rect 3850 2950 3950 3050
rect 3598 2878 3620 2912
rect 3654 2878 3678 2912
rect 3598 2840 3678 2878
rect 3800 2850 4000 2950
rect 4098 2912 4178 2958
rect 4098 2878 4120 2912
rect 4154 2878 4178 2912
rect 3598 2806 3620 2840
rect 3654 2806 3678 2840
rect 3598 2768 3678 2806
rect 3598 2734 3620 2768
rect 3654 2734 3678 2768
rect 3850 2750 3950 2850
rect 4098 2840 4178 2878
rect 4098 2806 4120 2840
rect 4154 2806 4178 2840
rect 4098 2768 4178 2806
rect 3598 2696 3678 2734
rect 3598 2662 3620 2696
rect 3654 2662 3678 2696
rect 3598 2624 3678 2662
rect 3800 2650 4000 2750
rect 4098 2734 4120 2768
rect 4154 2734 4178 2768
rect 4098 2696 4178 2734
rect 4098 2662 4120 2696
rect 4154 2662 4178 2696
rect 3598 2590 3620 2624
rect 3654 2590 3678 2624
rect 3598 2552 3678 2590
rect 3598 2518 3620 2552
rect 3654 2518 3678 2552
rect 3850 2550 3950 2650
rect 4098 2624 4178 2662
rect 4098 2590 4120 2624
rect 4154 2590 4178 2624
rect 4098 2552 4178 2590
rect 3598 2480 3678 2518
rect 3598 2446 3620 2480
rect 3654 2446 3678 2480
rect 3800 2450 4000 2550
rect 4098 2518 4120 2552
rect 4154 2518 4178 2552
rect 4098 2480 4178 2518
rect 3598 2408 3678 2446
rect 3598 2374 3620 2408
rect 3654 2374 3678 2408
rect 3598 2336 3678 2374
rect 3850 2350 3950 2450
rect 4098 2446 4120 2480
rect 4154 2446 4178 2480
rect 4098 2408 4178 2446
rect 4098 2374 4120 2408
rect 4154 2374 4178 2408
rect 3598 2302 3620 2336
rect 3654 2302 3678 2336
rect 3598 2264 3678 2302
rect 3598 2230 3620 2264
rect 3654 2230 3678 2264
rect 3800 2250 4000 2350
rect 4098 2336 4178 2374
rect 4098 2302 4120 2336
rect 4154 2302 4178 2336
rect 4098 2264 4178 2302
rect 3598 2192 3678 2230
rect 3598 2158 3620 2192
rect 3654 2158 3678 2192
rect 3598 2120 3678 2158
rect 3850 2150 3950 2250
rect 4098 2230 4120 2264
rect 4154 2230 4178 2264
rect 4098 2192 4178 2230
rect 4098 2158 4120 2192
rect 4154 2158 4178 2192
rect 3598 2086 3620 2120
rect 3654 2086 3678 2120
rect 3598 2040 3678 2086
rect 3800 2050 4000 2150
rect 4098 2120 4178 2158
rect 4098 2086 4120 2120
rect 4154 2086 4178 2120
rect 3850 1950 3950 2050
rect 4098 2040 4178 2086
rect 8422 2912 8502 2958
rect 8650 2950 8750 3050
rect 8422 2878 8444 2912
rect 8478 2878 8502 2912
rect 8422 2840 8502 2878
rect 8600 2850 8800 2950
rect 8922 2912 9002 2958
rect 8922 2878 8944 2912
rect 8978 2878 9002 2912
rect 8422 2806 8444 2840
rect 8478 2806 8502 2840
rect 8422 2768 8502 2806
rect 8422 2734 8444 2768
rect 8478 2734 8502 2768
rect 8650 2750 8750 2850
rect 8922 2840 9002 2878
rect 8922 2806 8944 2840
rect 8978 2806 9002 2840
rect 8922 2768 9002 2806
rect 8422 2696 8502 2734
rect 8422 2662 8444 2696
rect 8478 2662 8502 2696
rect 8422 2624 8502 2662
rect 8600 2650 8800 2750
rect 8922 2734 8944 2768
rect 8978 2734 9002 2768
rect 8922 2696 9002 2734
rect 8922 2662 8944 2696
rect 8978 2662 9002 2696
rect 8422 2590 8444 2624
rect 8478 2590 8502 2624
rect 8422 2552 8502 2590
rect 8422 2518 8444 2552
rect 8478 2518 8502 2552
rect 8650 2550 8750 2650
rect 8922 2624 9002 2662
rect 8922 2590 8944 2624
rect 8978 2590 9002 2624
rect 8922 2552 9002 2590
rect 8422 2480 8502 2518
rect 8422 2446 8444 2480
rect 8478 2446 8502 2480
rect 8600 2450 8800 2550
rect 8922 2518 8944 2552
rect 8978 2518 9002 2552
rect 8922 2480 9002 2518
rect 8422 2408 8502 2446
rect 8422 2374 8444 2408
rect 8478 2374 8502 2408
rect 8422 2336 8502 2374
rect 8650 2350 8750 2450
rect 8922 2446 8944 2480
rect 8978 2446 9002 2480
rect 8922 2408 9002 2446
rect 8922 2374 8944 2408
rect 8978 2374 9002 2408
rect 8422 2302 8444 2336
rect 8478 2302 8502 2336
rect 8422 2264 8502 2302
rect 8422 2230 8444 2264
rect 8478 2230 8502 2264
rect 8600 2250 8800 2350
rect 8922 2336 9002 2374
rect 8922 2302 8944 2336
rect 8978 2302 9002 2336
rect 8922 2264 9002 2302
rect 8422 2192 8502 2230
rect 8422 2158 8444 2192
rect 8478 2158 8502 2192
rect 8422 2120 8502 2158
rect 8650 2150 8750 2250
rect 8922 2230 8944 2264
rect 8978 2230 9002 2264
rect 8922 2192 9002 2230
rect 8922 2158 8944 2192
rect 8978 2158 9002 2192
rect 8422 2086 8444 2120
rect 8478 2086 8502 2120
rect 8422 2040 8502 2086
rect 8600 2050 8800 2150
rect 8922 2120 9002 2158
rect 8922 2086 8944 2120
rect 8978 2086 9002 2120
rect 8650 1950 8750 2050
rect 8922 2040 9002 2086
rect 11196 2912 11278 2958
rect 11450 2950 11550 3050
rect 11650 2950 11750 3050
rect 11850 2950 11950 3050
rect 12050 2950 12150 3050
rect 12250 2950 12350 3050
rect 12450 2950 12550 3050
rect 11196 2878 11220 2912
rect 11254 2878 11278 2912
rect 11196 2840 11278 2878
rect 11400 2850 12600 2950
rect 11196 2806 11220 2840
rect 11254 2806 11278 2840
rect 11196 2768 11278 2806
rect 11196 2734 11220 2768
rect 11254 2734 11278 2768
rect 11450 2750 11550 2850
rect 11650 2750 11750 2850
rect 11850 2750 11950 2850
rect 12050 2750 12150 2850
rect 12250 2750 12350 2850
rect 12450 2750 12550 2850
rect 11196 2696 11278 2734
rect 11196 2662 11220 2696
rect 11254 2662 11278 2696
rect 11196 2624 11278 2662
rect 11400 2650 12600 2750
rect 11196 2590 11220 2624
rect 11254 2590 11278 2624
rect 11196 2552 11278 2590
rect 11196 2518 11220 2552
rect 11254 2518 11278 2552
rect 11450 2550 11550 2650
rect 11650 2550 11750 2650
rect 11850 2550 11950 2650
rect 12050 2550 12150 2650
rect 12250 2550 12350 2650
rect 12450 2550 12550 2650
rect 11196 2480 11278 2518
rect 11196 2446 11220 2480
rect 11254 2446 11278 2480
rect 11400 2450 12600 2550
rect 11196 2408 11278 2446
rect 11196 2374 11220 2408
rect 11254 2374 11278 2408
rect 11196 2336 11278 2374
rect 11450 2350 11550 2450
rect 11650 2350 11750 2450
rect 11850 2350 11950 2450
rect 12050 2350 12150 2450
rect 12250 2350 12350 2450
rect 12450 2350 12550 2450
rect 11196 2302 11220 2336
rect 11254 2302 11278 2336
rect 11196 2264 11278 2302
rect 11196 2230 11220 2264
rect 11254 2230 11278 2264
rect 11400 2250 12600 2350
rect 11196 2192 11278 2230
rect 11196 2158 11220 2192
rect 11254 2158 11278 2192
rect 11196 2120 11278 2158
rect 11450 2150 11550 2250
rect 11650 2150 11750 2250
rect 11850 2150 11950 2250
rect 12050 2150 12150 2250
rect 12250 2150 12350 2250
rect 12450 2150 12550 2250
rect 11196 2086 11220 2120
rect 11254 2086 11278 2120
rect 11196 2040 11278 2086
rect 11400 2050 12600 2150
rect 11450 1950 11550 2050
rect 11650 1950 11750 2050
rect 11850 1950 11950 2050
rect 12050 1950 12150 2050
rect 12250 1950 12350 2050
rect 12450 1950 12550 2050
rect -200 1850 1200 1950
rect 3800 1850 4000 1950
rect 8600 1850 8800 1950
rect 11400 1850 12600 1950
rect -150 1750 -50 1850
rect 50 1750 150 1850
rect 250 1750 350 1850
rect 450 1750 550 1850
rect 650 1750 750 1850
rect 850 1750 950 1850
rect 1050 1750 1150 1850
rect 1250 1750 1350 1800
rect 1450 1750 1550 1800
rect 1650 1750 1750 1800
rect 1850 1750 1950 1800
rect 2050 1750 2150 1800
rect 2250 1750 2350 1800
rect 2450 1750 2550 1800
rect 2650 1750 2750 1800
rect 2850 1750 2950 1800
rect 3050 1750 3150 1800
rect 3250 1750 3350 1800
rect 3450 1750 3550 1800
rect 3650 1750 3750 1800
rect 3850 1750 3950 1850
rect 4050 1750 4150 1800
rect 4250 1750 4350 1800
rect 4450 1750 4550 1800
rect 4650 1750 4750 1800
rect 4850 1750 4950 1800
rect 5050 1750 5150 1800
rect 5250 1750 5350 1800
rect 5450 1750 5550 1800
rect 5650 1750 5750 1800
rect 5850 1750 5950 1800
rect 6050 1750 6150 1800
rect 6250 1750 6350 1800
rect 6450 1750 6550 1800
rect 6650 1750 6750 1800
rect 6850 1750 6950 1800
rect 7050 1750 7150 1800
rect 7250 1750 7350 1800
rect 7450 1750 7550 1800
rect 7650 1750 7750 1800
rect 7850 1750 7950 1800
rect 8050 1750 8150 1800
rect 8250 1750 8350 1800
rect 8450 1750 8550 1800
rect 8650 1750 8750 1850
rect 8850 1750 8950 1800
rect 9050 1750 9150 1800
rect 9250 1750 9350 1800
rect 9450 1750 9550 1800
rect 9650 1750 9750 1800
rect 9850 1750 9950 1800
rect 10050 1750 10150 1800
rect 10250 1750 10350 1800
rect 10450 1750 10550 1800
rect 10650 1750 10750 1800
rect 10850 1750 10950 1800
rect 11050 1750 11150 1800
rect 11250 1750 11350 1800
rect 11450 1750 11550 1850
rect 11650 1750 11750 1850
rect 11850 1750 11950 1850
rect 12050 1750 12150 1850
rect 12250 1750 12350 1850
rect 12450 1750 12550 1850
rect -200 1650 12600 1750
rect -150 1550 -50 1650
rect 50 1550 150 1650
rect 250 1600 350 1650
rect 450 1600 550 1650
rect 650 1600 750 1650
rect 850 1600 950 1650
rect 1050 1600 1150 1650
rect 1250 1600 1350 1650
rect 1450 1600 1550 1650
rect 1650 1600 1750 1650
rect 1850 1600 1950 1650
rect 2050 1600 2150 1650
rect 2250 1600 2350 1650
rect 2450 1600 2550 1650
rect 2650 1600 2750 1650
rect 2850 1600 2950 1650
rect 3050 1600 3150 1650
rect 3250 1600 3350 1650
rect 3450 1600 3550 1650
rect 3650 1600 3750 1650
rect 3850 1600 3950 1650
rect 4050 1600 4150 1650
rect 4250 1600 4350 1650
rect 4450 1600 4550 1650
rect 4650 1600 4750 1650
rect 4850 1600 4950 1650
rect 5050 1600 5150 1650
rect 5250 1600 5350 1650
rect 5450 1600 5550 1650
rect 5650 1600 5750 1650
rect 5850 1600 5950 1650
rect 6050 1550 6150 1650
rect 6250 1550 6350 1650
rect 6450 1600 6550 1650
rect 6650 1600 6750 1650
rect 6850 1600 6950 1650
rect 7050 1600 7150 1650
rect 7250 1600 7350 1650
rect 7450 1600 7550 1650
rect 7650 1600 7750 1650
rect 7850 1600 7950 1650
rect 8050 1600 8150 1650
rect 8250 1600 8350 1650
rect 8450 1600 8550 1650
rect 8650 1600 8750 1650
rect 8850 1600 8950 1650
rect 9050 1600 9150 1650
rect 9250 1600 9350 1650
rect 9450 1600 9550 1650
rect 9650 1600 9750 1650
rect 9850 1600 9950 1650
rect 10050 1600 10150 1650
rect 10250 1600 10350 1650
rect 10450 1600 10550 1650
rect 10650 1600 10750 1650
rect 10850 1600 10950 1650
rect 11050 1600 11150 1650
rect 11250 1600 11350 1650
rect 11450 1600 11550 1650
rect 11650 1600 11750 1650
rect 11850 1600 11950 1650
rect 12050 1600 12150 1650
rect 12250 1550 12350 1650
rect 12450 1550 12550 1650
rect -200 1450 200 1550
rect 6000 1450 6400 1550
rect 12200 1450 12600 1550
rect -150 1350 -50 1450
rect 50 1350 150 1450
rect 386 1350 466 1364
rect -200 1312 466 1350
rect -200 1278 408 1312
rect 442 1278 466 1312
rect -200 1250 466 1278
rect -150 1150 -50 1250
rect 50 1150 150 1250
rect 386 1240 466 1250
rect 386 1206 408 1240
rect 442 1206 466 1240
rect 386 1168 466 1206
rect 386 1150 408 1168
rect -200 1134 408 1150
rect 442 1134 466 1168
rect -200 1096 466 1134
rect -200 1062 408 1096
rect 442 1062 466 1096
rect -200 1050 466 1062
rect -150 950 -50 1050
rect 50 950 150 1050
rect 386 1024 466 1050
rect 386 990 408 1024
rect 442 990 466 1024
rect 386 952 466 990
rect 386 950 408 952
rect -200 918 408 950
rect 442 918 466 952
rect -200 880 466 918
rect -200 850 408 880
rect -150 750 -50 850
rect 50 750 150 850
rect 386 846 408 850
rect 442 846 466 880
rect 386 808 466 846
rect 386 774 408 808
rect 442 774 466 808
rect 386 750 466 774
rect -200 736 466 750
rect -200 702 408 736
rect 442 702 466 736
rect -200 664 466 702
rect -200 650 408 664
rect -150 550 -50 650
rect 50 550 150 650
rect 386 630 408 650
rect 442 630 466 664
rect 386 592 466 630
rect 386 558 408 592
rect 442 558 466 592
rect 386 550 466 558
rect -200 520 466 550
rect -200 486 408 520
rect 442 486 466 520
rect -200 450 466 486
rect -150 350 -50 450
rect 50 350 150 450
rect 386 436 466 450
rect 5734 1350 5814 1364
rect 6050 1350 6150 1450
rect 6250 1350 6350 1450
rect 6586 1350 6666 1364
rect 5734 1312 6666 1350
rect 5734 1278 5756 1312
rect 5790 1278 6608 1312
rect 6642 1278 6666 1312
rect 5734 1250 6666 1278
rect 5734 1240 5814 1250
rect 5734 1206 5756 1240
rect 5790 1206 5814 1240
rect 5734 1168 5814 1206
rect 5734 1134 5756 1168
rect 5790 1150 5814 1168
rect 6050 1150 6150 1250
rect 6250 1150 6350 1250
rect 6586 1240 6666 1250
rect 6586 1206 6608 1240
rect 6642 1206 6666 1240
rect 6586 1168 6666 1206
rect 6586 1150 6608 1168
rect 5790 1134 6608 1150
rect 6642 1134 6666 1168
rect 5734 1096 6666 1134
rect 5734 1062 5756 1096
rect 5790 1062 6608 1096
rect 6642 1062 6666 1096
rect 5734 1050 6666 1062
rect 5734 1024 5814 1050
rect 5734 990 5756 1024
rect 5790 990 5814 1024
rect 5734 952 5814 990
rect 5734 918 5756 952
rect 5790 950 5814 952
rect 6050 950 6150 1050
rect 6250 950 6350 1050
rect 6586 1024 6666 1050
rect 6586 990 6608 1024
rect 6642 990 6666 1024
rect 6586 952 6666 990
rect 6586 950 6608 952
rect 5790 918 6608 950
rect 6642 918 6666 952
rect 5734 880 6666 918
rect 5734 846 5756 880
rect 5790 850 6608 880
rect 5790 846 5814 850
rect 5734 808 5814 846
rect 5734 774 5756 808
rect 5790 774 5814 808
rect 5734 750 5814 774
rect 6050 750 6150 850
rect 6250 750 6350 850
rect 6586 846 6608 850
rect 6642 846 6666 880
rect 6586 808 6666 846
rect 6586 774 6608 808
rect 6642 774 6666 808
rect 6586 750 6666 774
rect 5734 736 6666 750
rect 5734 702 5756 736
rect 5790 702 6608 736
rect 6642 702 6666 736
rect 5734 664 6666 702
rect 5734 630 5756 664
rect 5790 650 6608 664
rect 5790 630 5814 650
rect 5734 592 5814 630
rect 5734 558 5756 592
rect 5790 558 5814 592
rect 5734 550 5814 558
rect 6050 550 6150 650
rect 6250 550 6350 650
rect 6586 630 6608 650
rect 6642 630 6666 664
rect 6586 592 6666 630
rect 6586 558 6608 592
rect 6642 558 6666 592
rect 6586 550 6666 558
rect 5734 520 6666 550
rect 5734 486 5756 520
rect 5790 486 6608 520
rect 6642 486 6666 520
rect 5734 450 6666 486
rect 5734 436 5814 450
rect 6050 350 6150 450
rect 6250 350 6350 450
rect 6586 436 6666 450
rect 11932 1350 12014 1364
rect 12250 1350 12350 1450
rect 12450 1350 12550 1450
rect 11932 1312 12600 1350
rect 11932 1278 11956 1312
rect 11990 1278 12600 1312
rect 11932 1250 12600 1278
rect 11932 1240 12014 1250
rect 11932 1206 11956 1240
rect 11990 1206 12014 1240
rect 11932 1168 12014 1206
rect 11932 1134 11956 1168
rect 11990 1150 12014 1168
rect 12250 1150 12350 1250
rect 12450 1150 12550 1250
rect 11990 1134 12600 1150
rect 11932 1096 12600 1134
rect 11932 1062 11956 1096
rect 11990 1062 12600 1096
rect 11932 1050 12600 1062
rect 11932 1024 12014 1050
rect 11932 990 11956 1024
rect 11990 990 12014 1024
rect 11932 952 12014 990
rect 11932 918 11956 952
rect 11990 950 12014 952
rect 12250 950 12350 1050
rect 12450 950 12550 1050
rect 11990 918 12600 950
rect 11932 880 12600 918
rect 11932 846 11956 880
rect 11990 850 12600 880
rect 11990 846 12014 850
rect 11932 808 12014 846
rect 11932 774 11956 808
rect 11990 774 12014 808
rect 11932 750 12014 774
rect 12250 750 12350 850
rect 12450 750 12550 850
rect 11932 736 12600 750
rect 11932 702 11956 736
rect 11990 702 12600 736
rect 11932 664 12600 702
rect 11932 630 11956 664
rect 11990 650 12600 664
rect 11990 630 12014 650
rect 11932 592 12014 630
rect 11932 558 11956 592
rect 11990 558 12014 592
rect 11932 550 12014 558
rect 12250 550 12350 650
rect 12450 550 12550 650
rect 11932 520 12600 550
rect 11932 486 11956 520
rect 11990 486 12600 520
rect 11932 450 12600 486
rect 11932 436 12014 450
rect 12250 350 12350 450
rect 12450 350 12550 450
rect -200 250 200 350
rect -150 150 -50 250
rect 50 150 150 250
rect 250 150 350 200
rect 450 150 550 200
rect 650 150 750 350
rect 850 150 950 350
rect 1050 150 1150 350
rect 1250 150 1350 350
rect 1450 150 1550 350
rect 1650 150 1750 350
rect 1850 150 1950 350
rect 2050 150 2150 350
rect 2250 150 2350 350
rect 2450 150 2550 350
rect 2650 150 2750 350
rect 2850 150 2950 350
rect 3050 150 3150 350
rect 3250 150 3350 350
rect 3450 150 3550 350
rect 3650 150 3750 350
rect 3850 150 3950 350
rect 4050 150 4150 350
rect 4250 150 4350 350
rect 4450 150 4550 350
rect 4650 150 4750 350
rect 4850 150 4950 350
rect 5050 150 5150 350
rect 5250 150 5350 350
rect 5450 150 5550 350
rect 6000 250 6400 350
rect 5650 150 5750 200
rect 5850 150 5950 200
rect 6050 150 6150 250
rect 6250 150 6350 250
rect 6450 150 6550 200
rect 6650 150 6750 200
rect 6850 150 6950 350
rect 7050 150 7150 350
rect 7250 150 7350 350
rect 7450 150 7550 350
rect 7650 150 7750 350
rect 7850 150 7950 350
rect 8050 150 8150 350
rect 8250 150 8350 350
rect 8450 150 8550 350
rect 8650 150 8750 350
rect 8850 150 8950 350
rect 9050 150 9150 350
rect 9250 150 9350 350
rect 9450 150 9550 350
rect 9650 150 9750 350
rect 9850 150 9950 350
rect 10050 150 10150 350
rect 10250 150 10350 350
rect 10450 150 10550 350
rect 10650 150 10750 350
rect 10850 150 10950 350
rect 11050 150 11150 350
rect 11250 150 11350 350
rect 11450 150 11550 350
rect 11650 150 11750 350
rect 12200 250 12600 350
rect 11850 150 11950 200
rect 12050 150 12150 200
rect 12250 150 12350 250
rect 12450 150 12550 250
rect -200 50 12600 150
rect -150 -50 -50 50
rect 50 -50 150 50
rect 250 -50 350 50
rect 450 -50 550 50
rect 650 -50 750 50
rect 850 -50 950 50
rect 1050 -50 1150 50
rect 1250 -50 1350 50
rect 1450 -50 1550 50
rect 1650 -50 1750 50
rect 1850 -50 1950 50
rect 2050 -50 2150 50
rect 2250 -50 2350 50
rect 2450 -50 2550 50
rect 2650 -50 2750 50
rect 2850 -50 2950 50
rect 3050 -50 3150 50
rect 3250 -50 3350 50
rect 3450 -50 3550 50
rect 3650 -50 3750 50
rect 3850 -50 3950 50
rect 4050 -50 4150 50
rect 4250 -50 4350 50
rect 4450 -50 4550 50
rect 4650 -50 4750 50
rect 4850 -50 4950 50
rect 5050 -50 5150 50
rect 5250 -50 5350 50
rect 5450 -50 5550 50
rect 5650 -50 5750 50
rect 5850 -50 5950 50
rect 6050 -50 6150 50
rect 6250 -50 6350 50
rect 6450 -50 6550 50
rect 6650 -50 6750 50
rect 6850 -50 6950 50
rect 7050 -50 7150 50
rect 7250 -50 7350 50
rect 7450 -50 7550 50
rect 7650 -50 7750 50
rect 7850 -50 7950 50
rect 8050 -50 8150 50
rect 8250 -50 8350 50
rect 8450 -50 8550 50
rect 8650 -50 8750 50
rect 8850 -50 8950 50
rect 9050 -50 9150 50
rect 9250 -50 9350 50
rect 9450 -50 9550 50
rect 9650 -50 9750 50
rect 9850 -50 9950 50
rect 10050 -50 10150 50
rect 10250 -50 10350 50
rect 10450 -50 10550 50
rect 10650 -50 10750 50
rect 10850 -50 10950 50
rect 11050 -50 11150 50
rect 11250 -50 11350 50
rect 11450 -50 11550 50
rect 11650 -50 11750 50
rect 11850 -50 11950 50
rect 12050 -50 12150 50
rect 12250 -50 12350 50
rect 12450 -50 12550 50
rect -200 -150 12600 -50
rect -150 -200 -50 -150
rect 50 -200 150 -150
rect 250 -200 350 -150
rect 450 -200 550 -150
rect 650 -200 750 -150
rect 850 -200 950 -150
rect 1050 -200 1150 -150
rect 1250 -200 1350 -150
rect 1450 -200 1550 -150
rect 1650 -200 1750 -150
rect 1850 -200 1950 -150
rect 2050 -200 2150 -150
rect 2250 -200 2350 -150
rect 2450 -200 2550 -150
rect 2650 -200 2750 -150
rect 2850 -200 2950 -150
rect 3050 -200 3150 -150
rect 3250 -200 3350 -150
rect 3450 -200 3550 -150
rect 3650 -200 3750 -150
rect 3850 -200 3950 -150
rect 4050 -200 4150 -150
rect 4250 -200 4350 -150
rect 4450 -200 4550 -150
rect 4650 -200 4750 -150
rect 4850 -200 4950 -150
rect 5050 -200 5150 -150
rect 5250 -200 5350 -150
rect 5450 -200 5550 -150
rect 5650 -200 5750 -150
rect 5850 -200 5950 -150
rect 6050 -200 6150 -150
rect 6250 -200 6350 -150
rect 6450 -200 6550 -150
rect 6650 -200 6750 -150
rect 6850 -200 6950 -150
rect 7050 -200 7150 -150
rect 7250 -200 7350 -150
rect 7450 -200 7550 -150
rect 7650 -200 7750 -150
rect 7850 -200 7950 -150
rect 8050 -200 8150 -150
rect 8250 -200 8350 -150
rect 8450 -200 8550 -150
rect 8650 -200 8750 -150
rect 8850 -200 8950 -150
rect 9050 -200 9150 -150
rect 9250 -200 9350 -150
rect 9450 -200 9550 -150
rect 9650 -200 9750 -150
rect 9850 -200 9950 -150
rect 10050 -200 10150 -150
rect 10250 -200 10350 -150
rect 10450 -200 10550 -150
rect 10650 -200 10750 -150
rect 10850 -200 10950 -150
rect 11050 -200 11150 -150
rect 11250 -200 11350 -150
rect 11450 -200 11550 -150
rect 11650 -200 11750 -150
rect 11850 -200 11950 -150
rect 12050 -200 12150 -150
rect 12250 -200 12350 -150
rect 12450 -200 12550 -150
<< metal2 >>
rect -150 3550 -50 3600
rect 50 3550 150 3600
rect 250 3550 350 3600
rect 450 3550 550 3600
rect 650 3550 750 3600
rect 850 3550 950 3600
rect 1050 3550 1150 3600
rect 1250 3550 1350 3600
rect 1450 3550 1550 3600
rect 1650 3550 1750 3600
rect 1850 3550 1950 3600
rect 2050 3550 2150 3600
rect 2250 3550 2350 3600
rect 2450 3550 2550 3600
rect 2650 3550 2750 3600
rect 2850 3550 2950 3600
rect 3050 3550 3150 3600
rect 3250 3550 3350 3600
rect 3450 3550 3550 3600
rect 3650 3550 3750 3600
rect 3850 3550 3950 3600
rect 4050 3550 4150 3600
rect 4250 3550 4350 3600
rect 4450 3550 4550 3600
rect 4650 3550 4750 3600
rect 4850 3550 4950 3600
rect 5050 3550 5150 3600
rect 5250 3550 5350 3600
rect 5450 3550 5550 3600
rect 5650 3550 5750 3600
rect 5850 3550 5950 3600
rect 6050 3550 6150 3600
rect 6250 3550 6350 3600
rect 6450 3550 6550 3600
rect 6650 3550 6750 3600
rect 6850 3550 6950 3600
rect 7050 3550 7150 3600
rect 7250 3550 7350 3600
rect 7450 3550 7550 3600
rect 7650 3550 7750 3600
rect 7850 3550 7950 3600
rect 8050 3550 8150 3600
rect 8250 3550 8350 3600
rect 8450 3550 8550 3600
rect 8650 3550 8750 3600
rect 8850 3550 8950 3600
rect 9050 3550 9150 3600
rect 9250 3550 9350 3600
rect 9450 3550 9550 3600
rect 9650 3550 9750 3600
rect 9850 3550 9950 3600
rect 10050 3550 10150 3600
rect 10250 3550 10350 3600
rect 10450 3550 10550 3600
rect 10650 3550 10750 3600
rect 10850 3550 10950 3600
rect 11050 3550 11150 3600
rect 11250 3550 11350 3600
rect 11450 3550 11550 3600
rect 11650 3550 11750 3600
rect 11850 3550 11950 3600
rect 12050 3550 12150 3600
rect 12250 3550 12350 3600
rect 12450 3550 12550 3600
rect -200 3450 12600 3550
rect -150 3350 -50 3450
rect 50 3350 150 3450
rect 250 3350 350 3450
rect 450 3350 550 3450
rect 650 3350 750 3450
rect 850 3350 950 3450
rect 1050 3350 1150 3450
rect 1250 3350 1350 3450
rect 1450 3350 1550 3450
rect 1650 3350 1750 3450
rect 1850 3350 1950 3450
rect 2050 3350 2150 3450
rect 2250 3350 2350 3450
rect 2450 3350 2550 3450
rect 2650 3350 2750 3450
rect 2850 3350 2950 3450
rect 3050 3350 3150 3450
rect 3250 3350 3350 3450
rect 3450 3350 3550 3450
rect 3650 3350 3750 3450
rect 3850 3350 3950 3450
rect 4050 3350 4150 3450
rect 4250 3350 4350 3450
rect 4450 3350 4550 3450
rect 4650 3350 4750 3450
rect 4850 3350 4950 3450
rect 5050 3350 5150 3450
rect 5250 3350 5350 3450
rect 5450 3350 5550 3450
rect 5650 3350 5750 3450
rect 5850 3350 5950 3450
rect 6050 3350 6150 3450
rect 6250 3350 6350 3450
rect 6450 3350 6550 3450
rect 6650 3350 6750 3450
rect 6850 3350 6950 3450
rect 7050 3350 7150 3450
rect 7250 3350 7350 3450
rect 7450 3350 7550 3450
rect 7650 3350 7750 3450
rect 7850 3350 7950 3450
rect 8050 3350 8150 3450
rect 8250 3350 8350 3450
rect 8450 3350 8550 3450
rect 8650 3350 8750 3450
rect 8850 3350 8950 3450
rect 9050 3350 9150 3450
rect 9250 3350 9350 3450
rect 9450 3350 9550 3450
rect 9650 3350 9750 3450
rect 9850 3350 9950 3450
rect 10050 3350 10150 3450
rect 10250 3350 10350 3450
rect 10450 3350 10550 3450
rect 10650 3350 10750 3450
rect 10850 3350 10950 3450
rect 11050 3350 11150 3450
rect 11250 3350 11350 3450
rect 11450 3350 11550 3450
rect 11650 3350 11750 3450
rect 11850 3350 11950 3450
rect 12050 3350 12150 3450
rect 12250 3350 12350 3450
rect 12450 3350 12550 3450
rect -200 3250 12600 3350
rect -150 3150 -50 3250
rect 50 3150 150 3250
rect 250 3150 350 3250
rect 450 3150 550 3250
rect 650 3150 750 3250
rect 850 3150 950 3250
rect 1050 3150 1150 3250
rect 1250 3200 1350 3250
rect 1450 3200 1550 3250
rect 1650 3200 1750 3250
rect 1850 3200 1950 3250
rect 2050 3200 2150 3250
rect 2250 3200 2350 3250
rect 2450 3200 2550 3250
rect 2650 3200 2750 3250
rect 2850 3200 2950 3250
rect 3050 3200 3150 3250
rect 3250 3200 3350 3250
rect 3450 3200 3550 3250
rect 3650 3200 3750 3250
rect 3850 3150 3950 3250
rect 4050 3200 4150 3250
rect 4250 3200 4350 3250
rect 4450 3200 4550 3250
rect 4650 3200 4750 3250
rect 4850 3200 4950 3250
rect 5050 3200 5150 3250
rect 5250 3200 5350 3250
rect 5450 3200 5550 3250
rect 5650 3200 5750 3250
rect 5850 3200 5950 3250
rect 6050 3200 6150 3250
rect 6250 3200 6350 3250
rect 6450 3200 6550 3250
rect 6650 3200 6750 3250
rect 6850 3200 6950 3250
rect 7050 3200 7150 3250
rect 7250 3200 7350 3250
rect 7450 3200 7550 3250
rect 7650 3200 7750 3250
rect 7850 3200 7950 3250
rect 8050 3200 8150 3250
rect 8250 3200 8350 3250
rect 8450 3200 8550 3250
rect 8650 3150 8750 3250
rect 8850 3200 8950 3250
rect 9050 3200 9150 3250
rect 9250 3200 9350 3250
rect 9450 3200 9550 3250
rect 9650 3200 9750 3250
rect 9850 3200 9950 3250
rect 10050 3200 10150 3250
rect 10250 3200 10350 3250
rect 10450 3200 10550 3250
rect 10650 3200 10750 3250
rect 10850 3200 10950 3250
rect 11050 3200 11150 3250
rect 11250 3200 11350 3250
rect 11450 3150 11550 3250
rect 11650 3150 11750 3250
rect 11850 3150 11950 3250
rect 12050 3150 12150 3250
rect 12250 3150 12350 3250
rect 12450 3150 12550 3250
rect -200 3050 1200 3150
rect 3800 3050 4000 3150
rect 8600 3050 8800 3150
rect 11400 3050 12600 3150
rect -150 2950 -50 3050
rect 50 2950 150 3050
rect 250 2950 350 3050
rect 450 2950 550 3050
rect 650 2950 750 3050
rect 850 2950 950 3050
rect 1050 2950 1150 3050
rect 1322 2950 1402 2958
rect -200 2850 1402 2950
rect 3598 2950 3678 2958
rect 3850 2950 3950 3050
rect 4098 2950 4178 2958
rect 2480 2880 2520 2920
rect -150 2750 -50 2850
rect 50 2750 150 2850
rect 250 2750 350 2850
rect 450 2750 550 2850
rect 650 2750 750 2850
rect 850 2750 950 2850
rect 1050 2750 1150 2850
rect 1322 2750 1402 2850
rect -200 2650 1402 2750
rect -150 2550 -50 2650
rect 50 2550 150 2650
rect 250 2550 350 2650
rect 450 2550 550 2650
rect 650 2550 750 2650
rect 850 2550 950 2650
rect 1050 2550 1150 2650
rect 1322 2550 1402 2650
rect -200 2450 1402 2550
rect -150 2350 -50 2450
rect 50 2350 150 2450
rect 250 2350 350 2450
rect 450 2350 550 2450
rect 650 2350 750 2450
rect 850 2350 950 2450
rect 1050 2350 1150 2450
rect 1322 2350 1402 2450
rect -200 2250 1402 2350
rect -150 2150 -50 2250
rect 50 2150 150 2250
rect 250 2150 350 2250
rect 450 2150 550 2250
rect 650 2150 750 2250
rect 850 2150 950 2250
rect 1050 2150 1150 2250
rect 1322 2150 1402 2250
rect -200 2050 1402 2150
rect -150 1950 -50 2050
rect 50 1950 150 2050
rect 250 1950 350 2050
rect 450 1950 550 2050
rect 650 1950 750 2050
rect 850 1950 950 2050
rect 1050 1950 1150 2050
rect 1322 2040 1402 2050
rect 3598 2850 4178 2950
rect 8422 2950 8502 2958
rect 8650 2950 8750 3050
rect 8922 2950 9002 2958
rect 6280 2880 6320 2920
rect 3598 2750 3678 2850
rect 3850 2750 3950 2850
rect 4098 2750 4178 2850
rect 3598 2650 4178 2750
rect 3598 2550 3678 2650
rect 3850 2550 3950 2650
rect 4098 2550 4178 2650
rect 3598 2450 4178 2550
rect 3598 2350 3678 2450
rect 3850 2350 3950 2450
rect 4098 2350 4178 2450
rect 3598 2250 4178 2350
rect 3598 2150 3678 2250
rect 3850 2150 3950 2250
rect 4098 2150 4178 2250
rect 3598 2050 4178 2150
rect 8422 2850 9002 2950
rect 11196 2950 11278 2958
rect 11450 2950 11550 3050
rect 11650 2950 11750 3050
rect 11850 2950 11950 3050
rect 12050 2950 12150 3050
rect 12250 2950 12350 3050
rect 12450 2950 12550 3050
rect 10080 2880 10120 2920
rect 8422 2750 8502 2850
rect 8650 2750 8750 2850
rect 8922 2750 9002 2850
rect 8422 2650 9002 2750
rect 8422 2550 8502 2650
rect 8650 2550 8750 2650
rect 8922 2550 9002 2650
rect 8422 2450 9002 2550
rect 8422 2350 8502 2450
rect 8650 2350 8750 2450
rect 8922 2350 9002 2450
rect 8422 2250 9002 2350
rect 8422 2150 8502 2250
rect 8650 2150 8750 2250
rect 8922 2150 9002 2250
rect 3598 2040 3678 2050
rect 3850 1950 3950 2050
rect 4098 2040 4178 2050
rect -200 1850 1200 1950
rect 3800 1850 4000 1950
rect -150 1750 -50 1850
rect 50 1750 150 1850
rect 250 1750 350 1850
rect 450 1750 550 1850
rect 650 1750 750 1850
rect 850 1750 950 1850
rect 1050 1750 1150 1850
rect 1250 1750 1350 1800
rect 1450 1750 1550 1800
rect 1650 1750 1750 1800
rect 1850 1750 1950 1800
rect 2050 1750 2150 1800
rect 2250 1750 2350 1800
rect 2450 1750 2550 1800
rect 2650 1750 2750 1800
rect 2850 1750 2950 1800
rect 3050 1750 3150 1800
rect 3250 1750 3350 1800
rect 3450 1750 3550 1800
rect 3650 1750 3750 1800
rect 3850 1750 3950 1850
rect 4050 1750 4150 1800
rect 4250 1750 4350 1800
rect 4450 1750 4550 2100
rect 4650 1750 4750 2100
rect 4850 1750 4950 2100
rect 5050 1750 5150 2100
rect 5250 1750 5350 2100
rect 5450 1750 5550 2100
rect 5650 1750 5750 2100
rect 5850 1750 5950 2100
rect 6050 1750 6150 2100
rect 6250 1750 6350 2100
rect 6450 1750 6550 2100
rect 6650 1750 6750 2100
rect 6850 1750 6950 2100
rect 7050 1750 7150 2100
rect 7250 1750 7350 2100
rect 7450 1750 7550 2100
rect 7650 1750 7750 2100
rect 7850 1750 7950 2100
rect 8050 1750 8150 2100
rect 8422 2050 9002 2150
rect 8422 2040 8502 2050
rect 8650 1950 8750 2050
rect 8922 2040 9002 2050
rect 11196 2850 12600 2950
rect 11196 2750 11278 2850
rect 11450 2750 11550 2850
rect 11650 2750 11750 2850
rect 11850 2750 11950 2850
rect 12050 2750 12150 2850
rect 12250 2750 12350 2850
rect 12450 2750 12550 2850
rect 11196 2650 12600 2750
rect 11196 2550 11278 2650
rect 11450 2550 11550 2650
rect 11650 2550 11750 2650
rect 11850 2550 11950 2650
rect 12050 2550 12150 2650
rect 12250 2550 12350 2650
rect 12450 2550 12550 2650
rect 11196 2450 12600 2550
rect 11196 2350 11278 2450
rect 11450 2350 11550 2450
rect 11650 2350 11750 2450
rect 11850 2350 11950 2450
rect 12050 2350 12150 2450
rect 12250 2350 12350 2450
rect 12450 2350 12550 2450
rect 11196 2250 12600 2350
rect 11196 2150 11278 2250
rect 11450 2150 11550 2250
rect 11650 2150 11750 2250
rect 11850 2150 11950 2250
rect 12050 2150 12150 2250
rect 12250 2150 12350 2250
rect 12450 2150 12550 2250
rect 11196 2050 12600 2150
rect 11196 2040 11278 2050
rect 11450 1950 11550 2050
rect 11650 1950 11750 2050
rect 11850 1950 11950 2050
rect 12050 1950 12150 2050
rect 12250 1950 12350 2050
rect 12450 1950 12550 2050
rect 8600 1850 8800 1950
rect 11400 1850 12600 1950
rect 8250 1750 8350 1800
rect 8450 1750 8550 1800
rect 8650 1750 8750 1850
rect 8850 1750 8950 1800
rect 9050 1750 9150 1800
rect 9250 1750 9350 1800
rect 9450 1750 9550 1800
rect 9650 1750 9750 1800
rect 9850 1750 9950 1800
rect 10050 1750 10150 1800
rect 10250 1750 10350 1800
rect 10450 1750 10550 1800
rect 10650 1750 10750 1800
rect 10850 1750 10950 1800
rect 11050 1750 11150 1800
rect 11250 1750 11350 1800
rect 11450 1750 11550 1850
rect 11650 1750 11750 1850
rect 11850 1750 11950 1850
rect 12050 1750 12150 1850
rect 12250 1750 12350 1850
rect 12450 1750 12550 1850
rect -200 1650 12600 1750
rect -150 1550 -50 1650
rect 50 1550 150 1650
rect 250 1600 350 1650
rect 450 1600 550 1650
rect 650 1600 750 1650
rect 850 1600 950 1650
rect 1050 1600 1150 1650
rect 1250 1600 1350 1650
rect 1450 1600 1550 1650
rect 1650 1600 1750 1650
rect 1850 1600 1950 1650
rect 2050 1600 2150 1650
rect 2250 1600 2350 1650
rect 2450 1600 2550 1650
rect 2650 1600 2750 1650
rect 2850 1600 2950 1650
rect 3050 1600 3150 1650
rect 3250 1600 3350 1650
rect 3450 1600 3550 1650
rect 3650 1600 3750 1650
rect 3850 1600 3950 1650
rect 4050 1600 4150 1650
rect 4250 1600 4350 1650
rect -200 1450 200 1550
rect 4450 1500 4550 1650
rect 4650 1500 4750 1650
rect 4850 1500 4950 1650
rect 5050 1500 5150 1650
rect 5250 1500 5350 1650
rect 5450 1500 5550 1650
rect 5650 1500 5750 1650
rect 5850 1500 5950 1650
rect 6050 1550 6150 1650
rect 6250 1550 6350 1650
rect 6000 1450 6400 1550
rect 6450 1500 6550 1650
rect 6650 1500 6750 1650
rect 6850 1500 6950 1650
rect 7050 1500 7150 1650
rect 7250 1500 7350 1650
rect 7450 1500 7550 1650
rect 7650 1500 7750 1650
rect 7850 1500 7950 1650
rect 8050 1500 8150 1650
rect 8250 1600 8350 1650
rect 8450 1600 8550 1650
rect 8650 1600 8750 1650
rect 8850 1600 8950 1650
rect 9050 1600 9150 1650
rect 9250 1600 9350 1650
rect 9450 1600 9550 1650
rect 9650 1600 9750 1650
rect 9850 1600 9950 1650
rect 10050 1600 10150 1650
rect 10250 1600 10350 1650
rect 10450 1600 10550 1650
rect 10650 1600 10750 1650
rect 10850 1600 10950 1650
rect 11050 1600 11150 1650
rect 11250 1600 11350 1650
rect 11450 1600 11550 1650
rect 11650 1600 11750 1650
rect 11850 1600 11950 1650
rect 12050 1600 12150 1650
rect 12250 1550 12350 1650
rect 12450 1550 12550 1650
rect 12200 1450 12600 1550
rect -150 1350 -50 1450
rect 50 1350 150 1450
rect 6050 1350 6150 1450
rect 6250 1350 6350 1450
rect 12250 1350 12350 1450
rect 12450 1350 12550 1450
rect -200 1250 200 1350
rect 6000 1250 6400 1350
rect 12200 1250 12600 1350
rect -150 1150 -50 1250
rect 50 1150 150 1250
rect 6050 1150 6150 1250
rect 6250 1150 6350 1250
rect 12250 1150 12350 1250
rect 12450 1150 12550 1250
rect -200 1050 200 1150
rect 6000 1050 6400 1150
rect 12200 1050 12600 1150
rect -150 950 -50 1050
rect 50 950 150 1050
rect 6050 950 6150 1050
rect 6250 950 6350 1050
rect 12250 950 12350 1050
rect 12450 950 12550 1050
rect -200 850 200 950
rect 6000 850 6400 950
rect 12200 850 12600 950
rect -150 750 -50 850
rect 50 750 150 850
rect 6050 750 6150 850
rect 6250 750 6350 850
rect 12250 750 12350 850
rect 12450 750 12550 850
rect -200 650 200 750
rect 6000 650 6400 750
rect 12200 650 12600 750
rect -150 550 -50 650
rect 50 550 150 650
rect 6050 550 6150 650
rect 6250 550 6350 650
rect 12250 550 12350 650
rect 12450 550 12550 650
rect -200 450 200 550
rect -150 350 -50 450
rect 50 350 150 450
rect -200 250 200 350
rect 650 300 750 500
rect 850 300 950 500
rect 1050 300 1150 500
rect 1250 300 1350 500
rect 1450 300 1550 500
rect 1650 300 1750 500
rect 1850 300 1950 500
rect 2050 300 2150 500
rect 2250 300 2350 500
rect 2450 300 2550 500
rect 2650 300 2750 500
rect 2850 300 2950 500
rect 3050 300 3150 500
rect 3250 300 3350 500
rect 3450 300 3550 500
rect 3650 300 3750 500
rect 3850 300 3950 500
rect 4050 300 4150 500
rect 4250 300 4350 500
rect 4450 300 4550 500
rect 4650 300 4750 500
rect 4850 300 4950 500
rect 5050 300 5150 500
rect 5250 300 5350 500
rect 5450 300 5550 500
rect 6000 450 6400 550
rect 6050 350 6150 450
rect 6250 350 6350 450
rect 6000 250 6400 350
rect 6850 300 6950 500
rect 7050 300 7150 500
rect 7250 300 7350 500
rect 7450 300 7550 500
rect 7650 300 7750 500
rect 7850 300 7950 500
rect 8050 300 8150 500
rect 8250 300 8350 500
rect 8450 300 8550 500
rect 8650 300 8750 500
rect 8850 300 8950 500
rect 9050 300 9150 500
rect 9250 300 9350 500
rect 9450 300 9550 500
rect 9650 300 9750 500
rect 9850 300 9950 500
rect 10050 300 10150 500
rect 10250 300 10350 500
rect 10450 300 10550 500
rect 10650 300 10750 500
rect 10850 300 10950 500
rect 11050 300 11150 500
rect 11250 300 11350 500
rect 11450 300 11550 500
rect 11650 300 11750 500
rect 12200 450 12600 550
rect 12250 350 12350 450
rect 12450 350 12550 450
rect 12200 250 12600 350
rect -150 150 -50 250
rect 50 150 150 250
rect 250 150 350 200
rect 450 150 550 200
rect 650 150 750 200
rect 850 150 950 200
rect 1050 150 1150 200
rect 1250 150 1350 200
rect 1450 150 1550 200
rect 1650 150 1750 200
rect 1850 150 1950 200
rect 2050 150 2150 200
rect 2250 150 2350 200
rect 2450 150 2550 200
rect 2650 150 2750 200
rect 2850 150 2950 200
rect 3050 150 3150 200
rect 3250 150 3350 200
rect 3450 150 3550 200
rect 3650 150 3750 200
rect 3850 150 3950 200
rect 4050 150 4150 200
rect 4250 150 4350 200
rect 4450 150 4550 200
rect 4650 150 4750 200
rect 4850 150 4950 200
rect 5050 150 5150 200
rect 5250 150 5350 200
rect 5450 150 5550 200
rect 5650 150 5750 200
rect 5850 150 5950 200
rect 6050 150 6150 250
rect 6250 150 6350 250
rect 6450 150 6550 200
rect 6650 150 6750 200
rect 6850 150 6950 200
rect 7050 150 7150 200
rect 7250 150 7350 200
rect 7450 150 7550 200
rect 7650 150 7750 200
rect 7850 150 7950 200
rect 8050 150 8150 200
rect 8250 150 8350 200
rect 8450 150 8550 200
rect 8650 150 8750 200
rect 8850 150 8950 200
rect 9050 150 9150 200
rect 9250 150 9350 200
rect 9450 150 9550 200
rect 9650 150 9750 200
rect 9850 150 9950 200
rect 10050 150 10150 200
rect 10250 150 10350 200
rect 10450 150 10550 200
rect 10650 150 10750 200
rect 10850 150 10950 200
rect 11050 150 11150 200
rect 11250 150 11350 200
rect 11450 150 11550 200
rect 11650 150 11750 200
rect 11850 150 11950 200
rect 12050 150 12150 200
rect 12250 150 12350 250
rect 12450 150 12550 250
rect -200 50 12600 150
rect -150 -50 -50 50
rect 50 -50 150 50
rect 250 -50 350 50
rect 450 -50 550 50
rect 650 -50 750 50
rect 850 -50 950 50
rect 1050 -50 1150 50
rect 1250 -50 1350 50
rect 1450 -50 1550 50
rect 1650 -50 1750 50
rect 1850 -50 1950 50
rect 2050 -50 2150 50
rect 2250 -50 2350 50
rect 2450 -50 2550 50
rect 2650 -50 2750 50
rect 2850 -50 2950 50
rect 3050 -50 3150 50
rect 3250 -50 3350 50
rect 3450 -50 3550 50
rect 3650 -50 3750 50
rect 3850 -50 3950 50
rect 4050 -50 4150 50
rect 4250 -50 4350 50
rect 4450 -50 4550 50
rect 4650 -50 4750 50
rect 4850 -50 4950 50
rect 5050 -50 5150 50
rect 5250 -50 5350 50
rect 5450 -50 5550 50
rect 5650 -50 5750 50
rect 5850 -50 5950 50
rect 6050 -50 6150 50
rect 6250 -50 6350 50
rect 6450 -50 6550 50
rect 6650 -50 6750 50
rect 6850 -50 6950 50
rect 7050 -50 7150 50
rect 7250 -50 7350 50
rect 7450 -50 7550 50
rect 7650 -50 7750 50
rect 7850 -50 7950 50
rect 8050 -50 8150 50
rect 8250 -50 8350 50
rect 8450 -50 8550 50
rect 8650 -50 8750 50
rect 8850 -50 8950 50
rect 9050 -50 9150 50
rect 9250 -50 9350 50
rect 9450 -50 9550 50
rect 9650 -50 9750 50
rect 9850 -50 9950 50
rect 10050 -50 10150 50
rect 10250 -50 10350 50
rect 10450 -50 10550 50
rect 10650 -50 10750 50
rect 10850 -50 10950 50
rect 11050 -50 11150 50
rect 11250 -50 11350 50
rect 11450 -50 11550 50
rect 11650 -50 11750 50
rect 11850 -50 11950 50
rect 12050 -50 12150 50
rect 12250 -50 12350 50
rect 12450 -50 12550 50
rect -200 -150 12600 -50
rect -150 -200 -50 -150
rect 50 -200 150 -150
rect 250 -200 350 -150
rect 450 -200 550 -150
rect 650 -200 750 -150
rect 850 -200 950 -150
rect 1050 -200 1150 -150
rect 1250 -200 1350 -150
rect 1450 -200 1550 -150
rect 1650 -200 1750 -150
rect 1850 -200 1950 -150
rect 2050 -200 2150 -150
rect 2250 -200 2350 -150
rect 2450 -200 2550 -150
rect 2650 -200 2750 -150
rect 2850 -200 2950 -150
rect 3050 -200 3150 -150
rect 3250 -200 3350 -150
rect 3450 -200 3550 -150
rect 3650 -200 3750 -150
rect 3850 -200 3950 -150
rect 4050 -200 4150 -150
rect 4250 -200 4350 -150
rect 4450 -200 4550 -150
rect 4650 -200 4750 -150
rect 4850 -200 4950 -150
rect 5050 -200 5150 -150
rect 5250 -200 5350 -150
rect 5450 -200 5550 -150
rect 5650 -200 5750 -150
rect 5850 -200 5950 -150
rect 6050 -200 6150 -150
rect 6250 -200 6350 -150
rect 6450 -200 6550 -150
rect 6650 -200 6750 -150
rect 6850 -200 6950 -150
rect 7050 -200 7150 -150
rect 7250 -200 7350 -150
rect 7450 -200 7550 -150
rect 7650 -200 7750 -150
rect 7850 -200 7950 -150
rect 8050 -200 8150 -150
rect 8250 -200 8350 -150
rect 8450 -200 8550 -150
rect 8650 -200 8750 -150
rect 8850 -200 8950 -150
rect 9050 -200 9150 -150
rect 9250 -200 9350 -150
rect 9450 -200 9550 -150
rect 9650 -200 9750 -150
rect 9850 -200 9950 -150
rect 10050 -200 10150 -150
rect 10250 -200 10350 -150
rect 10450 -200 10550 -150
rect 10650 -200 10750 -150
rect 10850 -200 10950 -150
rect 11050 -200 11150 -150
rect 11250 -200 11350 -150
rect 11450 -200 11550 -150
rect 11650 -200 11750 -150
rect 11850 -200 11950 -150
rect 12050 -200 12150 -150
rect 12250 -200 12350 -150
rect 12450 -200 12550 -150
<< metal3 >>
rect 2450 2450 2550 2550
rect 4250 2540 4350 2550
rect 3260 2460 4350 2540
rect 2460 1350 2540 2450
rect 3260 2150 3340 2460
rect 4250 2450 4350 2460
rect 8250 2540 8350 2550
rect 8250 2460 9340 2540
rect 8250 2450 8350 2460
rect 9260 2150 9340 2460
rect 10050 2450 10150 2550
rect 3250 2050 3350 2150
rect 9250 2050 9350 2150
rect 2450 1250 2550 1350
rect 3050 1250 3150 1350
rect 5450 1340 5550 1350
rect 6850 1340 6950 1350
rect 5450 1260 6950 1340
rect 5450 1250 5550 1260
rect 6850 1250 6950 1260
rect 3060 950 3140 1250
rect 10060 950 10140 2450
rect 3050 850 3150 950
rect 10050 850 10150 950
use via_M1_M2_1_a  NoName_294
timestamp 1508605124
transform 1 0 1362 0 1 2500
box -32 -32 32 32
use via_M1_M2_1_b  NoName_295
timestamp 1508605124
transform 1 0 1362 0 1 2628
box -32 -32 32 32
use via_M1_M2_1_c  NoName_296
timestamp 1508605124
transform 1 0 1362 0 1 2372
box -32 -32 32 32
use via_M1_M2_1_d  NoName_297
timestamp 1508605124
transform 1 0 1362 0 1 2756
box -32 -32 32 32
use via_M1_M2_1_e  NoName_298
timestamp 1508605124
transform 1 0 1362 0 1 2244
box -32 -32 32 32
use via_M1_M2_1_f  NoName_299
timestamp 1508605124
transform 1 0 1362 0 1 2884
box -32 -32 32 32
use via_M1_M2_1_g  NoName_300
timestamp 1508605124
transform 1 0 1362 0 1 2116
box -32 -32 32 32
use via_M1_M2_1_h  NoName_301
timestamp 1508605124
transform 1 0 3638 0 1 2500
box -32 -32 32 32
use via_M1_M2_1_i  NoName_302
timestamp 1508605124
transform 1 0 3638 0 1 2628
box -32 -32 32 32
use via_M1_M2_1_j  NoName_303
timestamp 1508605124
transform 1 0 3638 0 1 2372
box -32 -32 32 32
use via_M1_M2_1_k  NoName_304
timestamp 1508605124
transform 1 0 3638 0 1 2756
box -32 -32 32 32
use via_M1_M2_1_l  NoName_305
timestamp 1508605124
transform 1 0 3638 0 1 2244
box -32 -32 32 32
use via_M1_M2_1_m  NoName_306
timestamp 1508605124
transform 1 0 3638 0 1 2884
box -32 -32 32 32
use via_M1_M2_1_n  NoName_307
timestamp 1508605124
transform 1 0 3638 0 1 2116
box -32 -32 32 32
use via_M1_M2_1_o  NoName_308
timestamp 1508605124
transform 1 0 8962 0 1 2500
box -32 -32 32 32
use via_M1_M2_1_p  NoName_309
timestamp 1508605124
transform 1 0 8962 0 1 2628
box -32 -32 32 32
use via_M1_M2_1_q  NoName_310
timestamp 1508605124
transform 1 0 8962 0 1 2372
box -32 -32 32 32
use via_M1_M2_1_r  NoName_311
timestamp 1508605124
transform 1 0 8962 0 1 2756
box -32 -32 32 32
use via_M1_M2_1_s  NoName_312
timestamp 1508605124
transform 1 0 8962 0 1 2244
box -32 -32 32 32
use via_M1_M2_1_t  NoName_313
timestamp 1508605124
transform 1 0 8962 0 1 2884
box -32 -32 32 32
use via_M1_M2_1_u  NoName_314
timestamp 1508605124
transform 1 0 8962 0 1 2116
box -32 -32 32 32
use via_M1_M2_1_v  NoName_315
timestamp 1508605124
transform 1 0 11238 0 1 2500
box -32 -32 32 32
use via_M1_M2_1_w  NoName_316
timestamp 1508605124
transform 1 0 11238 0 1 2628
box -32 -32 32 32
use via_M1_M2_1_x  NoName_317
timestamp 1508605124
transform 1 0 11238 0 1 2372
box -32 -32 32 32
use via_M1_M2_1_y  NoName_318
timestamp 1508605124
transform 1 0 11238 0 1 2756
box -32 -32 32 32
use via_M1_M2_1_z  NoName_319
timestamp 1508605124
transform 1 0 11238 0 1 2244
box -32 -32 32 32
use via_M1_M2_1_{  NoName_320
timestamp 1508605124
transform 1 0 11238 0 1 2884
box -32 -32 32 32
use via_M1_M2_1_|  NoName_321
timestamp 1508605124
transform 1 0 11238 0 1 2116
box -32 -32 32 32
use via_M1_M2_1_}  NoName_322
timestamp 1508605124
transform 1 0 4138 0 1 2500
box -32 -32 32 32
use via_M1_M2_1_~  NoName_323
timestamp 1508605124
transform 1 0 4138 0 1 2628
box -32 -32 32 32
use XXXXX88  NoName_324
timestamp 1508605124
transform 1 0 4138 0 1 2372
box -32 -32 32 32
use XXXXX87  NoName_325
timestamp 1508605124
transform 1 0 4138 0 1 2756
box -32 -32 32 32
use XXXXX64  NoName_326
timestamp 1508605124
transform 1 0 4138 0 1 2244
box -32 -32 32 32
use XXXXX86  NoName_327
timestamp 1508605124
transform 1 0 4138 0 1 2884
box -32 -32 32 32
use XXXXX65  NoName_328
timestamp 1508605124
transform 1 0 4138 0 1 2116
box -32 -32 32 32
use XXXXX91  NoName_329
timestamp 1508605124
transform 1 0 8462 0 1 2500
box -32 -32 32 32
use XXXXX92  NoName_330
timestamp 1508605124
transform 1 0 8462 0 1 2628
box -32 -32 32 32
use XXXXX93  NoName_331
timestamp 1508605124
transform 1 0 8462 0 1 2372
box -32 -32 32 32
use XXXXX94  NoName_332
timestamp 1508605124
transform 1 0 8462 0 1 2756
box -32 -32 32 32
use XXXXX69  NoName_333
timestamp 1508605124
transform 1 0 8462 0 1 2244
box -32 -32 32 32
use XXXXX95  NoName_334
timestamp 1508605124
transform 1 0 8462 0 1 2884
box -32 -32 32 32
use XXXXX68  NoName_335
timestamp 1508605124
transform 1 0 8462 0 1 2116
box -32 -32 32 32
use via_M2_M3_0  NoName_336
timestamp 1508605124
transform 1 0 10100 0 1 2500
box -38 -38 38 38
use via_M2_M3_0  NoName_337
timestamp 1508605124
transform 1 0 10100 0 1 900
box -38 -38 38 38
use via_M2_M3_0  NoName_340
timestamp 1508605124
transform 1 0 3100 0 1 900
box -38 -38 38 38
use via_M2_M3_0  NoName_341
timestamp 1508605124
transform 1 0 3100 0 1 1300
box -38 -38 38 38
use via_M2_M3_0  NoName_344
timestamp 1508605124
transform 1 0 2500 0 1 2500
box -38 -38 38 38
use via_M2_M3_0  NoName_345
timestamp 1508605124
transform 1 0 2500 0 1 1300
box -38 -38 38 38
use via_M2_M3_0  NoName_348
timestamp 1508605124
transform 1 0 5500 0 1 1300
box -38 -38 38 38
use via_M2_M3_0  NoName_349
timestamp 1508605124
transform 1 0 6900 0 1 1300
box -38 -38 38 38
use via_M2_M3_0  NoName_352
timestamp 1508605124
transform 1 0 3300 0 1 2100
box -38 -38 38 38
use via_M2_M3_0  NoName_353
timestamp 1508605124
transform 1 0 4300 0 1 2500
box -38 -38 38 38
use via_M2_M3_0  NoName_356
timestamp 1508605124
transform 1 0 9300 0 1 2100
box -38 -38 38 38
use via_M2_M3_0  NoName_357
timestamp 1508605124
transform 1 0 8300 0 1 2500
box -38 -38 38 38
use XXXXX2  NoName_360
timestamp 1508605124
transform 1 0 700 0 1 350
box -32 -32 32 32
use XXXXX3  NoName_361
timestamp 1508605124
transform 1 0 900 0 1 350
box -32 -32 32 32
use XXXXX4  NoName_362
timestamp 1508605124
transform 1 0 1100 0 1 350
box -32 -32 32 32
use XXXXX5  NoName_363
timestamp 1508605124
transform 1 0 1300 0 1 350
box -32 -32 32 32
use XXXXX7  NoName_364
timestamp 1508605124
transform 1 0 1500 0 1 350
box -32 -32 32 32
use XXXXX6  NoName_365
timestamp 1508605124
transform 1 0 1700 0 1 350
box -32 -32 32 32
use XXXXX8  NoName_366
timestamp 1508605124
transform 1 0 1900 0 1 350
box -32 -32 32 32
use XXXXX9  NoName_367
timestamp 1508605124
transform 1 0 2100 0 1 350
box -32 -32 32 32
use XXXXX10  NoName_368
timestamp 1508605124
transform 1 0 2300 0 1 350
box -32 -32 32 32
use XXXXX11  NoName_369
timestamp 1508605124
transform 1 0 2500 0 1 350
box -32 -32 32 32
use XXXXX12  NoName_370
timestamp 1508605124
transform 1 0 2700 0 1 350
box -32 -32 32 32
use XXXXX13  NoName_371
timestamp 1508605124
transform 1 0 2900 0 1 350
box -32 -32 32 32
use XXXXX14  NoName_372
timestamp 1508605124
transform 1 0 3100 0 1 350
box -32 -32 32 32
use XXXXX15  NoName_373
timestamp 1508605124
transform 1 0 3300 0 1 350
box -32 -32 32 32
use XXXXX16  NoName_374
timestamp 1508605124
transform 1 0 3500 0 1 350
box -32 -32 32 32
use XXXXX17  NoName_375
timestamp 1508605124
transform 1 0 3700 0 1 350
box -32 -32 32 32
use XXXXX19  NoName_376
timestamp 1508605124
transform 1 0 3900 0 1 350
box -32 -32 32 32
use XXXXX18  NoName_377
timestamp 1508605124
transform 1 0 4100 0 1 350
box -32 -32 32 32
use XXXXX20  NoName_378
timestamp 1508605124
transform 1 0 4300 0 1 350
box -32 -32 32 32
use XXXXX21  NoName_379
timestamp 1508605124
transform 1 0 4500 0 1 350
box -32 -32 32 32
use XXXXX22  NoName_380
timestamp 1508605124
transform 1 0 4700 0 1 350
box -32 -32 32 32
use XXXXX23  NoName_381
timestamp 1508605124
transform 1 0 4900 0 1 350
box -32 -32 32 32
use XXXXX24  NoName_382
timestamp 1508605124
transform 1 0 5100 0 1 350
box -32 -32 32 32
use XXXXX25  NoName_383
timestamp 1508605124
transform 1 0 5300 0 1 350
box -32 -32 32 32
use XXXXX26  NoName_384
timestamp 1508605124
transform 1 0 5500 0 1 350
box -32 -32 32 32
use XXXXX31  NoName_385
timestamp 1508605124
transform 1 0 6900 0 1 350
box -32 -32 32 32
use XXXXX32  NoName_386
timestamp 1508605124
transform 1 0 7100 0 1 350
box -32 -32 32 32
use XXXXX34  NoName_387
timestamp 1508605124
transform 1 0 7300 0 1 350
box -32 -32 32 32
use XXXXX33  NoName_388
timestamp 1508605124
transform 1 0 7500 0 1 350
box -32 -32 32 32
use XXXXX35  NoName_389
timestamp 1508605124
transform 1 0 7700 0 1 350
box -32 -32 32 32
use XXXXX36  NoName_390
timestamp 1508605124
transform 1 0 7900 0 1 350
box -32 -32 32 32
use XXXXX37  NoName_391
timestamp 1508605124
transform 1 0 8100 0 1 350
box -32 -32 32 32
use XXXXX38  NoName_392
timestamp 1508605124
transform 1 0 8300 0 1 350
box -32 -32 32 32
use XXXXX39  NoName_393
timestamp 1508605124
transform 1 0 8500 0 1 350
box -32 -32 32 32
use XXXXX41  NoName_394
timestamp 1508605124
transform 1 0 8700 0 1 350
box -32 -32 32 32
use XXXXX40  NoName_395
timestamp 1508605124
transform 1 0 8900 0 1 350
box -32 -32 32 32
use XXXXX42  NoName_396
timestamp 1508605124
transform 1 0 9100 0 1 350
box -32 -32 32 32
use XXXXX43  NoName_397
timestamp 1508605124
transform 1 0 9300 0 1 350
box -32 -32 32 32
use XXXXX44  NoName_398
timestamp 1508605124
transform 1 0 9500 0 1 350
box -32 -32 32 32
use XXXXX45  NoName_399
timestamp 1508605124
transform 1 0 9700 0 1 350
box -32 -32 32 32
use XXXXX47  NoName_400
timestamp 1508605124
transform 1 0 9900 0 1 350
box -32 -32 32 32
use XXXXX46  NoName_401
timestamp 1508605124
transform 1 0 10100 0 1 350
box -32 -32 32 32
use XXXXX48  NoName_402
timestamp 1508605124
transform 1 0 10300 0 1 350
box -32 -32 32 32
use XXXXX49  NoName_403
timestamp 1508605124
transform 1 0 10500 0 1 350
box -32 -32 32 32
use XXXXX50  NoName_404
timestamp 1508605124
transform 1 0 10700 0 1 350
box -32 -32 32 32
use XXXXX51  NoName_405
timestamp 1508605124
transform 1 0 10900 0 1 350
box -32 -32 32 32
use XXXXX53  NoName_406
timestamp 1508605124
transform 1 0 11100 0 1 350
box -32 -32 32 32
use XXXXX52  NoName_407
timestamp 1508605124
transform 1 0 11300 0 1 350
box -32 -32 32 32
use XXXXX57  NoName_408
timestamp 1508605124
transform 1 0 11500 0 1 350
box -32 -32 32 32
use XXXXX56  NoName_409
timestamp 1508605124
transform 1 0 11700 0 1 350
box -32 -32 32 32
use XM1  XM1
timestamp 1508605124
transform 1 0 2500 0 1 2500
box -1181 -519 1181 519
use XM2  XM2
timestamp 1508605124
transform 1 0 3100 0 1 900
box -2727 -534 2727 534
use XM3  XM3
timestamp 1508605124
transform 1 0 10100 0 1 2500
box -1181 -519 1181 519
use XM4  XM4
timestamp 1508605124
transform 1 0 9300 0 1 900
box -2727 -534 2727 534
use XM5  XM5
timestamp 1508605124
transform 1 0 6300 0 1 2500
box -2205 -519 2205 519
<< labels >>
flabel metal3 s 10100 1700 10100 1700 0 FreeSans 2000 0 0 0 out
port 1 nsew
flabel metal2 s 2480 2880 2520 2920 0 FreeSans 2000 0 0 0 ia
port 2 nsew
flabel metal2 s 10080 2880 10120 2920 0 FreeSans 2000 0 0 0 ib
port 3 nsew
flabel metal2 s 6280 2880 6320 2920 0 FreeSans 2000 0 0 0 icmbias
port 4 nsew
flabel metal2 s 3100 500 3100 500 0 FreeSans 2000 0 0 0 vdd
port 5 nsew
flabel metal2 s 9300 500 9300 500 0 FreeSans 2000 0 0 0 vdd
port 5 nsew
flabel metal2 s 6300 2100 6300 2100 0 FreeSans 2000 0 0 0 vss
port 6 nsew
<< end >>
