magic
tech sky130A
magscale 1 2
timestamp 1679988683
<< checkpaint >>
rect -2451 -1789 2451 1789
<< pwell >>
rect -1191 -529 1191 529
<< nmoslvt >>
rect -995 -381 -925 319
rect -867 -381 -797 319
rect -739 -381 -669 319
rect -611 -381 -541 319
rect -483 -381 -413 319
rect -355 -381 -285 319
rect -227 -381 -157 319
rect -99 -381 -29 319
rect 29 -381 99 319
rect 157 -381 227 319
rect 285 -381 355 319
rect 413 -381 483 319
rect 541 -381 611 319
rect 669 -381 739 319
rect 797 -381 867 319
rect 925 -381 995 319
<< ndiff >>
rect -1053 307 -995 319
rect -1053 -369 -1041 307
rect -1007 -369 -995 307
rect -1053 -381 -995 -369
rect -925 307 -867 319
rect -925 -369 -913 307
rect -879 -369 -867 307
rect -925 -381 -867 -369
rect -797 307 -739 319
rect -797 -369 -785 307
rect -751 -369 -739 307
rect -797 -381 -739 -369
rect -669 307 -611 319
rect -669 -369 -657 307
rect -623 -369 -611 307
rect -669 -381 -611 -369
rect -541 307 -483 319
rect -541 -369 -529 307
rect -495 -369 -483 307
rect -541 -381 -483 -369
rect -413 307 -355 319
rect -413 -369 -401 307
rect -367 -369 -355 307
rect -413 -381 -355 -369
rect -285 307 -227 319
rect -285 -369 -273 307
rect -239 -369 -227 307
rect -285 -381 -227 -369
rect -157 307 -99 319
rect -157 -369 -145 307
rect -111 -369 -99 307
rect -157 -381 -99 -369
rect -29 307 29 319
rect -29 -369 -17 307
rect 17 -369 29 307
rect -29 -381 29 -369
rect 99 307 157 319
rect 99 -369 111 307
rect 145 -369 157 307
rect 99 -381 157 -369
rect 227 307 285 319
rect 227 -369 239 307
rect 273 -369 285 307
rect 227 -381 285 -369
rect 355 307 413 319
rect 355 -369 367 307
rect 401 -369 413 307
rect 355 -381 413 -369
rect 483 307 541 319
rect 483 -369 495 307
rect 529 -369 541 307
rect 483 -381 541 -369
rect 611 307 669 319
rect 611 -369 623 307
rect 657 -369 669 307
rect 611 -381 669 -369
rect 739 307 797 319
rect 739 -369 751 307
rect 785 -369 797 307
rect 739 -381 797 -369
rect 867 307 925 319
rect 867 -369 879 307
rect 913 -369 925 307
rect 867 -381 925 -369
rect 995 307 1053 319
rect 995 -369 1007 307
rect 1041 -369 1053 307
rect 995 -381 1053 -369
<< ndiffc >>
rect -1041 -369 -1007 307
rect -913 -369 -879 307
rect -785 -369 -751 307
rect -657 -369 -623 307
rect -529 -369 -495 307
rect -401 -369 -367 307
rect -273 -369 -239 307
rect -145 -369 -111 307
rect -17 -369 17 307
rect 111 -369 145 307
rect 239 -369 273 307
rect 367 -369 401 307
rect 495 -369 529 307
rect 623 -369 657 307
rect 751 -369 785 307
rect 879 -369 913 307
rect 1007 -369 1041 307
<< psubdiff >>
rect -1155 459 -1059 493
rect 1059 459 1155 493
rect -1155 397 -1121 459
rect 1121 397 1155 459
rect -1155 -459 -1121 -397
rect 1121 -459 1155 -397
rect -1155 -493 -1059 -459
rect 1059 -493 1155 -459
<< psubdiffcont >>
rect -1059 459 1059 493
rect -1155 -397 -1121 397
rect 1121 -397 1155 397
rect -1059 -493 1059 -459
<< poly >>
rect -995 391 -925 407
rect -995 357 -979 391
rect -941 357 -925 391
rect -995 319 -925 357
rect -867 391 -797 407
rect -867 357 -851 391
rect -813 357 -797 391
rect -867 319 -797 357
rect -739 391 -669 407
rect -739 357 -723 391
rect -685 357 -669 391
rect -739 319 -669 357
rect -611 391 -541 407
rect -611 357 -595 391
rect -557 357 -541 391
rect -611 319 -541 357
rect -483 391 -413 407
rect -483 357 -467 391
rect -429 357 -413 391
rect -483 319 -413 357
rect -355 391 -285 407
rect -355 357 -339 391
rect -301 357 -285 391
rect -355 319 -285 357
rect -227 391 -157 407
rect -227 357 -211 391
rect -173 357 -157 391
rect -227 319 -157 357
rect -99 391 -29 407
rect -99 357 -83 391
rect -45 357 -29 391
rect -99 319 -29 357
rect 29 391 99 407
rect 29 357 45 391
rect 83 357 99 391
rect 29 319 99 357
rect 157 391 227 407
rect 157 357 173 391
rect 211 357 227 391
rect 157 319 227 357
rect 285 391 355 407
rect 285 357 301 391
rect 339 357 355 391
rect 285 319 355 357
rect 413 391 483 407
rect 413 357 429 391
rect 467 357 483 391
rect 413 319 483 357
rect 541 391 611 407
rect 541 357 557 391
rect 595 357 611 391
rect 541 319 611 357
rect 669 391 739 407
rect 669 357 685 391
rect 723 357 739 391
rect 669 319 739 357
rect 797 391 867 407
rect 797 357 813 391
rect 851 357 867 391
rect 797 319 867 357
rect 925 391 995 407
rect 925 357 941 391
rect 979 357 995 391
rect 925 319 995 357
rect -995 -407 -925 -381
rect -867 -407 -797 -381
rect -739 -407 -669 -381
rect -611 -407 -541 -381
rect -483 -407 -413 -381
rect -355 -407 -285 -381
rect -227 -407 -157 -381
rect -99 -407 -29 -381
rect 29 -407 99 -381
rect 157 -407 227 -381
rect 285 -407 355 -381
rect 413 -407 483 -381
rect 541 -407 611 -381
rect 669 -407 739 -381
rect 797 -407 867 -381
rect 925 -407 995 -381
<< polycont >>
rect -979 357 -941 391
rect -851 357 -813 391
rect -723 357 -685 391
rect -595 357 -557 391
rect -467 357 -429 391
rect -339 357 -301 391
rect -211 357 -173 391
rect -83 357 -45 391
rect 45 357 83 391
rect 173 357 211 391
rect 301 357 339 391
rect 429 357 467 391
rect 557 357 595 391
rect 685 357 723 391
rect 813 357 851 391
rect 941 357 979 391
<< locali >>
rect -1155 459 -1059 493
rect 1059 459 1155 493
rect -1155 397 -1121 459
rect 1121 397 1155 459
rect -995 357 -979 391
rect -941 357 -925 391
rect -867 357 -851 391
rect -813 357 -797 391
rect -739 357 -723 391
rect -685 357 -669 391
rect -611 357 -595 391
rect -557 357 -541 391
rect -483 357 -467 391
rect -429 357 -413 391
rect -355 357 -339 391
rect -301 357 -285 391
rect -227 357 -211 391
rect -173 357 -157 391
rect -99 357 -83 391
rect -45 357 -29 391
rect 29 357 45 391
rect 83 357 99 391
rect 157 357 173 391
rect 211 357 227 391
rect 285 357 301 391
rect 339 357 355 391
rect 413 357 429 391
rect 467 357 483 391
rect 541 357 557 391
rect 595 357 611 391
rect 669 357 685 391
rect 723 357 739 391
rect 797 357 813 391
rect 851 357 867 391
rect 925 357 941 391
rect 979 357 995 391
rect -1041 307 -1007 323
rect -1041 -385 -1007 -369
rect -913 307 -879 323
rect -913 -385 -879 -369
rect -785 307 -751 323
rect -785 -385 -751 -369
rect -657 307 -623 323
rect -657 -385 -623 -369
rect -529 307 -495 323
rect -529 -385 -495 -369
rect -401 307 -367 323
rect -401 -385 -367 -369
rect -273 307 -239 323
rect -273 -385 -239 -369
rect -145 307 -111 323
rect -145 -385 -111 -369
rect -17 307 17 323
rect -17 -385 17 -369
rect 111 307 145 323
rect 111 -385 145 -369
rect 239 307 273 323
rect 239 -385 273 -369
rect 367 307 401 323
rect 367 -385 401 -369
rect 495 307 529 323
rect 495 -385 529 -369
rect 623 307 657 323
rect 623 -385 657 -369
rect 751 307 785 323
rect 751 -385 785 -369
rect 879 307 913 323
rect 879 -385 913 -369
rect 1007 307 1041 323
rect 1007 -385 1041 -369
rect -1155 -459 -1121 -397
rect 1121 -459 1155 -397
rect -1155 -493 -1059 -459
rect 1059 -493 1155 -459
<< viali >>
rect -979 357 -941 391
rect -851 357 -813 391
rect -723 357 -685 391
rect -595 357 -557 391
rect -467 357 -429 391
rect -339 357 -301 391
rect -211 357 -173 391
rect -83 357 -45 391
rect 45 357 83 391
rect 173 357 211 391
rect 301 357 339 391
rect 429 357 467 391
rect 557 357 595 391
rect 685 357 723 391
rect 813 357 851 391
rect 941 357 979 391
rect -1041 -369 -1007 307
rect -913 -369 -879 307
rect -785 -369 -751 307
rect -657 -369 -623 307
rect -529 -369 -495 307
rect -401 -369 -367 307
rect -273 -369 -239 307
rect -145 -369 -111 307
rect -17 -369 17 307
rect 111 -369 145 307
rect 239 -369 273 307
rect 367 -369 401 307
rect 495 -369 529 307
rect 623 -369 657 307
rect 751 -369 785 307
rect 879 -369 913 307
rect 1007 -369 1041 307
<< metal1 >>
rect -991 391 -929 397
rect -991 357 -979 391
rect -941 357 -929 391
rect -991 351 -929 357
rect -863 391 -801 397
rect -863 357 -851 391
rect -813 357 -801 391
rect -863 351 -801 357
rect -735 391 -673 397
rect -735 357 -723 391
rect -685 357 -673 391
rect -735 351 -673 357
rect -607 391 -545 397
rect -607 357 -595 391
rect -557 357 -545 391
rect -607 351 -545 357
rect -479 391 -417 397
rect -479 357 -467 391
rect -429 357 -417 391
rect -479 351 -417 357
rect -351 391 -289 397
rect -351 357 -339 391
rect -301 357 -289 391
rect -351 351 -289 357
rect -223 391 -161 397
rect -223 357 -211 391
rect -173 357 -161 391
rect -223 351 -161 357
rect -95 391 -33 397
rect -95 357 -83 391
rect -45 357 -33 391
rect -95 351 -33 357
rect 33 391 95 397
rect 33 357 45 391
rect 83 357 95 391
rect 33 351 95 357
rect 161 391 223 397
rect 161 357 173 391
rect 211 357 223 391
rect 161 351 223 357
rect 289 391 351 397
rect 289 357 301 391
rect 339 357 351 391
rect 289 351 351 357
rect 417 391 479 397
rect 417 357 429 391
rect 467 357 479 391
rect 417 351 479 357
rect 545 391 607 397
rect 545 357 557 391
rect 595 357 607 391
rect 545 351 607 357
rect 673 391 735 397
rect 673 357 685 391
rect 723 357 735 391
rect 673 351 735 357
rect 801 391 863 397
rect 801 357 813 391
rect 851 357 863 391
rect 801 351 863 357
rect 929 391 991 397
rect 929 357 941 391
rect 979 357 991 391
rect 929 351 991 357
rect -1047 307 -1001 319
rect -1047 -369 -1041 307
rect -1007 -369 -1001 307
rect -1047 -381 -1001 -369
rect -919 307 -873 319
rect -919 -369 -913 307
rect -879 -369 -873 307
rect -919 -381 -873 -369
rect -791 307 -745 319
rect -791 -369 -785 307
rect -751 -369 -745 307
rect -791 -381 -745 -369
rect -663 307 -617 319
rect -663 -369 -657 307
rect -623 -369 -617 307
rect -663 -381 -617 -369
rect -535 307 -489 319
rect -535 -369 -529 307
rect -495 -369 -489 307
rect -535 -381 -489 -369
rect -407 307 -361 319
rect -407 -369 -401 307
rect -367 -369 -361 307
rect -407 -381 -361 -369
rect -279 307 -233 319
rect -279 -369 -273 307
rect -239 -369 -233 307
rect -279 -381 -233 -369
rect -151 307 -105 319
rect -151 -369 -145 307
rect -111 -369 -105 307
rect -151 -381 -105 -369
rect -23 307 23 319
rect -23 -369 -17 307
rect 17 -369 23 307
rect -23 -381 23 -369
rect 105 307 151 319
rect 105 -369 111 307
rect 145 -369 151 307
rect 105 -381 151 -369
rect 233 307 279 319
rect 233 -369 239 307
rect 273 -369 279 307
rect 233 -381 279 -369
rect 361 307 407 319
rect 361 -369 367 307
rect 401 -369 407 307
rect 361 -381 407 -369
rect 489 307 535 319
rect 489 -369 495 307
rect 529 -369 535 307
rect 489 -381 535 -369
rect 617 307 663 319
rect 617 -369 623 307
rect 657 -369 663 307
rect 617 -381 663 -369
rect 745 307 791 319
rect 745 -369 751 307
rect 785 -369 791 307
rect 745 -381 791 -369
rect 873 307 919 319
rect 873 -369 879 307
rect 913 -369 919 307
rect 873 -381 919 -369
rect 1001 307 1047 319
rect 1001 -369 1007 307
rect 1041 -369 1047 307
rect 1001 -381 1047 -369
<< labels >>
flabel metal1 -960 374 -960 374 0 FreeSans 240 0 0 0 G
flabel metal1 -832 374 -832 374 0 FreeSans 240 0 0 0 G
flabel metal1 -704 374 -704 374 0 FreeSans 240 0 0 0 G
flabel metal1 -576 374 -576 374 0 FreeSans 240 0 0 0 G
flabel metal1 -448 374 -448 374 0 FreeSans 240 0 0 0 G
flabel metal1 -320 374 -320 374 0 FreeSans 240 0 0 0 G
flabel metal1 -192 374 -192 374 0 FreeSans 240 0 0 0 G
flabel metal1 -64 374 -64 374 0 FreeSans 240 0 0 0 G
flabel metal1 64 374 64 374 0 FreeSans 240 0 0 0 G
flabel metal1 192 374 192 374 0 FreeSans 240 0 0 0 G
flabel metal1 320 374 320 374 0 FreeSans 240 0 0 0 G
flabel metal1 448 374 448 374 0 FreeSans 240 0 0 0 G
flabel metal1 576 374 576 374 0 FreeSans 240 0 0 0 G
flabel metal1 704 374 704 374 0 FreeSans 240 0 0 0 G
flabel metal1 832 374 832 374 0 FreeSans 240 0 0 0 G
flabel metal1 960 374 960 374 0 FreeSans 240 0 0 0 G
flabel metal1 -1024 -31 -1024 -31 0 FreeSans 240 0 0 0 D
flabel metal1 -896 -31 -896 -31 0 FreeSans 240 0 0 0 S
flabel metal1 -768 -31 -768 -31 0 FreeSans 240 0 0 0 D
flabel metal1 -640 -31 -640 -31 0 FreeSans 240 0 0 0 S
flabel metal1 -512 -31 -512 -31 0 FreeSans 240 0 0 0 D
flabel metal1 -384 -31 -384 -31 0 FreeSans 240 0 0 0 S
flabel metal1 -256 -31 -256 -31 0 FreeSans 240 0 0 0 D
flabel metal1 -128 -31 -128 -31 0 FreeSans 240 0 0 0 S
flabel metal1 0 -31 0 -31 0 FreeSans 240 0 0 0 D
flabel metal1 128 -31 128 -31 0 FreeSans 240 0 0 0 S
flabel metal1 256 -31 256 -31 0 FreeSans 240 0 0 0 D
flabel metal1 384 -31 384 -31 0 FreeSans 240 0 0 0 S
flabel metal1 512 -31 512 -31 0 FreeSans 240 0 0 0 D
flabel metal1 640 -31 640 -31 0 FreeSans 240 0 0 0 S
flabel metal1 768 -31 768 -31 0 FreeSans 240 0 0 0 D
flabel metal1 896 -31 896 -31 0 FreeSans 240 0 0 0 S
flabel metal1 1024 -31 1024 -31 0 FreeSans 240 0 0 0 D
<< properties >>
string FIXED_BBOX -1138 -476 1138 476
<< end >>

