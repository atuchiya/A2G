magic
tech sky130A
magscale 1 2
timestamp 1679394724
<< checkpaint >>
rect -1210 4610 15010 4660
rect -1260 -1210 15060 4610
rect -1260 -1260 15010 -1210
<< viali >>
rect 344 2878 378 2912
rect 2620 2878 2654 2912
rect 4720 2878 4754 2912
rect 9044 2878 9078 2912
rect 11144 2878 11178 2912
rect 13420 2878 13454 2912
rect 344 2806 378 2840
rect 2620 2806 2654 2840
rect 4720 2806 4754 2840
rect 9044 2806 9078 2840
rect 11144 2806 11178 2840
rect 13420 2806 13454 2840
rect 344 2734 378 2768
rect 2620 2734 2654 2768
rect 4720 2734 4754 2768
rect 9044 2734 9078 2768
rect 11144 2734 11178 2768
rect 13420 2734 13454 2768
rect 344 2662 378 2696
rect 2620 2662 2654 2696
rect 4720 2662 4754 2696
rect 9044 2662 9078 2696
rect 11144 2662 11178 2696
rect 13420 2662 13454 2696
rect 344 2590 378 2624
rect 2620 2590 2654 2624
rect 4720 2590 4754 2624
rect 9044 2590 9078 2624
rect 11144 2590 11178 2624
rect 13420 2590 13454 2624
rect 344 2518 378 2552
rect 2620 2518 2654 2552
rect 4720 2518 4754 2552
rect 9044 2518 9078 2552
rect 11144 2518 11178 2552
rect 13420 2518 13454 2552
rect 344 2446 378 2480
rect 2620 2446 2654 2480
rect 4720 2446 4754 2480
rect 9044 2446 9078 2480
rect 11144 2446 11178 2480
rect 13420 2446 13454 2480
rect 344 2374 378 2408
rect 2620 2374 2654 2408
rect 4720 2374 4754 2408
rect 9044 2374 9078 2408
rect 11144 2374 11178 2408
rect 13420 2374 13454 2408
rect 344 2302 378 2336
rect 2620 2302 2654 2336
rect 4720 2302 4754 2336
rect 9044 2302 9078 2336
rect 11144 2302 11178 2336
rect 13420 2302 13454 2336
rect 344 2230 378 2264
rect 2620 2230 2654 2264
rect 4720 2230 4754 2264
rect 9044 2230 9078 2264
rect 11144 2230 11178 2264
rect 13420 2230 13454 2264
rect 344 2158 378 2192
rect 2620 2158 2654 2192
rect 4720 2158 4754 2192
rect 9044 2158 9078 2192
rect 11144 2158 11178 2192
rect 13420 2158 13454 2192
rect 344 2086 378 2120
rect 2620 2086 2654 2120
rect 4720 2086 4754 2120
rect 9044 2086 9078 2120
rect 11144 2086 11178 2120
rect 13420 2086 13454 2120
rect 1008 1278 1042 1312
rect 6356 1278 6390 1312
rect 7408 1278 7442 1312
rect 12756 1278 12790 1312
rect 1008 1206 1042 1240
rect 6356 1206 6390 1240
rect 7408 1206 7442 1240
rect 12756 1206 12790 1240
rect 1008 1134 1042 1168
rect 6356 1134 6390 1168
rect 7408 1134 7442 1168
rect 12756 1134 12790 1168
rect 1008 1062 1042 1096
rect 6356 1062 6390 1096
rect 7408 1062 7442 1096
rect 12756 1062 12790 1096
rect 1008 990 1042 1024
rect 6356 990 6390 1024
rect 7408 990 7442 1024
rect 12756 990 12790 1024
rect 1008 918 1042 952
rect 6356 918 6390 952
rect 7408 918 7442 952
rect 12756 918 12790 952
rect 1008 846 1042 880
rect 6356 846 6390 880
rect 7408 846 7442 880
rect 12756 846 12790 880
rect 1008 774 1042 808
rect 6356 774 6390 808
rect 7408 774 7442 808
rect 12756 774 12790 808
rect 1008 702 1042 736
rect 6356 702 6390 736
rect 7408 702 7442 736
rect 12756 702 12790 736
rect 1008 630 1042 664
rect 6356 630 6390 664
rect 7408 630 7442 664
rect 12756 630 12790 664
rect 1008 558 1042 592
rect 6356 558 6390 592
rect 7408 558 7442 592
rect 12756 558 12790 592
rect 1008 486 1042 520
rect 6356 486 6390 520
rect 7408 486 7442 520
rect 12756 486 12790 520
<< metal1 >>
rect 50 3350 150 3400
rect 250 3350 350 3400
rect 450 3350 550 3400
rect 650 3350 750 3400
rect 850 3350 950 3400
rect 1050 3350 1150 3400
rect 1250 3350 1350 3400
rect 1450 3350 1550 3400
rect 1650 3350 1750 3400
rect 1850 3350 1950 3400
rect 2050 3350 2150 3400
rect 2250 3350 2350 3400
rect 2450 3350 2550 3400
rect 2650 3350 2750 3400
rect 2850 3350 2950 3400
rect 3050 3350 3150 3400
rect 3250 3350 3350 3400
rect 3450 3350 3550 3400
rect 3650 3350 3750 3400
rect 3850 3350 3950 3400
rect 4050 3350 4150 3400
rect 4250 3350 4350 3400
rect 4450 3350 4550 3400
rect 4650 3350 4750 3400
rect 4850 3350 4950 3400
rect 5050 3350 5150 3400
rect 5250 3350 5350 3400
rect 5450 3350 5550 3400
rect 5650 3350 5750 3400
rect 5850 3350 5950 3400
rect 6050 3350 6150 3400
rect 6250 3350 6350 3400
rect 6450 3350 6550 3400
rect 6650 3350 6750 3400
rect 6850 3350 6950 3400
rect 7050 3350 7150 3400
rect 7250 3350 7350 3400
rect 7450 3350 7550 3400
rect 7650 3350 7750 3400
rect 7850 3350 7950 3400
rect 8050 3350 8150 3400
rect 8250 3350 8350 3400
rect 8450 3350 8550 3400
rect 8650 3350 8750 3400
rect 8850 3350 8950 3400
rect 9050 3350 9150 3400
rect 9250 3350 9350 3400
rect 9450 3350 9550 3400
rect 9650 3350 9750 3400
rect 9850 3350 9950 3400
rect 10050 3350 10150 3400
rect 10250 3350 10350 3400
rect 10450 3350 10550 3400
rect 10650 3350 10750 3400
rect 10850 3350 10950 3400
rect 11050 3350 11150 3400
rect 11250 3350 11350 3400
rect 11450 3350 11550 3400
rect 11650 3350 11750 3400
rect 11850 3350 11950 3400
rect 12050 3350 12150 3400
rect 12250 3350 12350 3400
rect 12450 3350 12550 3400
rect 12650 3350 12750 3400
rect 12850 3350 12950 3400
rect 13050 3350 13150 3400
rect 13250 3350 13350 3400
rect 13450 3350 13550 3400
rect 13650 3350 13750 3400
rect 0 3250 13800 3350
rect 50 3150 150 3250
rect 250 3150 350 3250
rect 450 3150 550 3250
rect 650 3150 750 3250
rect 850 3150 950 3250
rect 1050 3150 1150 3250
rect 1250 3150 1350 3250
rect 1450 3150 1550 3250
rect 1650 3150 1750 3250
rect 1850 3150 1950 3250
rect 2050 3150 2150 3250
rect 2250 3150 2350 3250
rect 2450 3150 2550 3250
rect 2650 3150 2750 3250
rect 2850 3150 2950 3250
rect 3050 3150 3150 3250
rect 3250 3150 3350 3250
rect 3450 3150 3550 3250
rect 3650 3150 3750 3250
rect 3850 3150 3950 3250
rect 4050 3150 4150 3250
rect 4250 3150 4350 3250
rect 4450 3150 4550 3250
rect 4650 3150 4750 3250
rect 4850 3150 4950 3250
rect 5050 3150 5150 3250
rect 5250 3150 5350 3250
rect 5450 3150 5550 3250
rect 5650 3150 5750 3250
rect 5850 3150 5950 3250
rect 6050 3150 6150 3250
rect 6250 3150 6350 3250
rect 6450 3150 6550 3250
rect 6650 3150 6750 3250
rect 6850 3150 6950 3250
rect 7050 3150 7150 3250
rect 7250 3150 7350 3250
rect 7450 3150 7550 3250
rect 7650 3150 7750 3250
rect 7850 3150 7950 3250
rect 8050 3150 8150 3250
rect 8250 3150 8350 3250
rect 8450 3150 8550 3250
rect 8650 3150 8750 3250
rect 8850 3150 8950 3250
rect 9050 3150 9150 3250
rect 9250 3150 9350 3250
rect 9450 3150 9550 3250
rect 9650 3150 9750 3250
rect 9850 3150 9950 3250
rect 10050 3150 10150 3250
rect 10250 3150 10350 3250
rect 10450 3150 10550 3250
rect 10650 3150 10750 3250
rect 10850 3150 10950 3250
rect 11050 3150 11150 3250
rect 11250 3150 11350 3250
rect 11450 3150 11550 3250
rect 11650 3150 11750 3250
rect 11850 3150 11950 3250
rect 12050 3150 12150 3250
rect 12250 3150 12350 3250
rect 12450 3150 12550 3250
rect 12650 3150 12750 3250
rect 12850 3150 12950 3250
rect 13050 3150 13150 3250
rect 13250 3150 13350 3250
rect 13450 3150 13550 3250
rect 13650 3150 13750 3250
rect 0 3050 13800 3150
rect 50 2950 150 3050
rect 0 2850 150 2950
rect 50 2750 150 2850
rect 0 2650 150 2750
rect 50 2550 150 2650
rect 0 2450 150 2550
rect 50 2350 150 2450
rect 0 2250 150 2350
rect 50 2150 150 2250
rect 0 2050 150 2150
rect 50 1950 150 2050
rect 320 2912 400 2958
rect 320 2878 344 2912
rect 378 2878 400 2912
rect 320 2840 400 2878
rect 320 2806 344 2840
rect 378 2806 400 2840
rect 320 2768 400 2806
rect 320 2734 344 2768
rect 378 2734 400 2768
rect 320 2696 400 2734
rect 320 2662 344 2696
rect 378 2662 400 2696
rect 320 2624 400 2662
rect 320 2590 344 2624
rect 378 2590 400 2624
rect 320 2552 400 2590
rect 320 2518 344 2552
rect 378 2518 400 2552
rect 320 2480 400 2518
rect 320 2446 344 2480
rect 378 2446 400 2480
rect 320 2408 400 2446
rect 320 2374 344 2408
rect 378 2374 400 2408
rect 320 2336 400 2374
rect 320 2302 344 2336
rect 378 2302 400 2336
rect 320 2264 400 2302
rect 320 2230 344 2264
rect 378 2230 400 2264
rect 320 2192 400 2230
rect 320 2158 344 2192
rect 378 2158 400 2192
rect 320 2120 400 2158
rect 320 2086 344 2120
rect 378 2086 400 2120
rect 320 2040 400 2086
rect 2598 2912 2678 2958
rect 2598 2878 2620 2912
rect 2654 2878 2678 2912
rect 2598 2840 2678 2878
rect 2598 2806 2620 2840
rect 2654 2806 2678 2840
rect 2598 2768 2678 2806
rect 2598 2734 2620 2768
rect 2654 2734 2678 2768
rect 2598 2696 2678 2734
rect 2598 2662 2620 2696
rect 2654 2662 2678 2696
rect 2598 2624 2678 2662
rect 2598 2590 2620 2624
rect 2654 2590 2678 2624
rect 2598 2552 2678 2590
rect 2598 2518 2620 2552
rect 2654 2518 2678 2552
rect 2598 2480 2678 2518
rect 2598 2446 2620 2480
rect 2654 2446 2678 2480
rect 2598 2408 2678 2446
rect 2598 2374 2620 2408
rect 2654 2374 2678 2408
rect 2598 2336 2678 2374
rect 2598 2302 2620 2336
rect 2654 2302 2678 2336
rect 2598 2264 2678 2302
rect 2598 2230 2620 2264
rect 2654 2230 2678 2264
rect 2598 2192 2678 2230
rect 2598 2158 2620 2192
rect 2654 2158 2678 2192
rect 2598 2120 2678 2158
rect 2598 2086 2620 2120
rect 2654 2086 2678 2120
rect 2598 2040 2678 2086
rect 2850 2950 2950 3050
rect 3050 2950 3150 3050
rect 3250 2950 3350 3050
rect 3450 2950 3550 3050
rect 3650 2950 3750 3050
rect 3850 2950 3950 3050
rect 4050 2950 4150 3050
rect 4250 2950 4350 3050
rect 4450 2950 4550 3050
rect 2850 2850 4550 2950
rect 2850 2750 2950 2850
rect 3050 2750 3150 2850
rect 3250 2750 3350 2850
rect 3450 2750 3550 2850
rect 3650 2750 3750 2850
rect 3850 2750 3950 2850
rect 4050 2750 4150 2850
rect 4250 2750 4350 2850
rect 4450 2750 4550 2850
rect 2850 2650 4550 2750
rect 2850 2550 2950 2650
rect 3050 2550 3150 2650
rect 3250 2550 3350 2650
rect 3450 2550 3550 2650
rect 3650 2550 3750 2650
rect 3850 2550 3950 2650
rect 4050 2550 4150 2650
rect 4250 2550 4350 2650
rect 4450 2550 4550 2650
rect 2850 2450 4550 2550
rect 2850 2350 2950 2450
rect 3050 2350 3150 2450
rect 3250 2350 3350 2450
rect 3450 2350 3550 2450
rect 3650 2350 3750 2450
rect 3850 2350 3950 2450
rect 4050 2350 4150 2450
rect 4250 2350 4350 2450
rect 4450 2350 4550 2450
rect 2850 2250 4550 2350
rect 2850 2150 2950 2250
rect 3050 2150 3150 2250
rect 3250 2150 3350 2250
rect 3450 2150 3550 2250
rect 3650 2150 3750 2250
rect 3850 2150 3950 2250
rect 4050 2150 4150 2250
rect 4250 2150 4350 2250
rect 4450 2150 4550 2250
rect 2850 2050 4550 2150
rect 2850 1950 2950 2050
rect 3050 1950 3150 2050
rect 3250 1950 3350 2050
rect 3450 1950 3550 2050
rect 3650 1950 3750 2050
rect 3850 1950 3950 2050
rect 4050 1950 4150 2050
rect 4250 1950 4350 2050
rect 4450 1950 4550 2050
rect 4698 2912 4778 2958
rect 4698 2878 4720 2912
rect 4754 2878 4778 2912
rect 4698 2840 4778 2878
rect 4698 2806 4720 2840
rect 4754 2806 4778 2840
rect 4698 2768 4778 2806
rect 4698 2734 4720 2768
rect 4754 2734 4778 2768
rect 4698 2696 4778 2734
rect 4698 2662 4720 2696
rect 4754 2662 4778 2696
rect 4698 2624 4778 2662
rect 4698 2590 4720 2624
rect 4754 2590 4778 2624
rect 4698 2552 4778 2590
rect 4698 2518 4720 2552
rect 4754 2518 4778 2552
rect 4698 2480 4778 2518
rect 4698 2446 4720 2480
rect 4754 2446 4778 2480
rect 4698 2408 4778 2446
rect 4698 2374 4720 2408
rect 4754 2374 4778 2408
rect 4698 2336 4778 2374
rect 4698 2302 4720 2336
rect 4754 2302 4778 2336
rect 4698 2264 4778 2302
rect 4698 2230 4720 2264
rect 4754 2230 4778 2264
rect 4698 2192 4778 2230
rect 4698 2158 4720 2192
rect 4754 2158 4778 2192
rect 4698 2120 4778 2158
rect 4698 2086 4720 2120
rect 4754 2086 4778 2120
rect 4698 2040 4778 2086
rect 9022 2912 9102 2958
rect 9022 2878 9044 2912
rect 9078 2878 9102 2912
rect 9022 2840 9102 2878
rect 9022 2806 9044 2840
rect 9078 2806 9102 2840
rect 9022 2768 9102 2806
rect 9022 2734 9044 2768
rect 9078 2734 9102 2768
rect 9022 2696 9102 2734
rect 9022 2662 9044 2696
rect 9078 2662 9102 2696
rect 9022 2624 9102 2662
rect 9022 2590 9044 2624
rect 9078 2590 9102 2624
rect 9022 2552 9102 2590
rect 9022 2518 9044 2552
rect 9078 2518 9102 2552
rect 9022 2480 9102 2518
rect 9022 2446 9044 2480
rect 9078 2446 9102 2480
rect 9022 2408 9102 2446
rect 9022 2374 9044 2408
rect 9078 2374 9102 2408
rect 9022 2336 9102 2374
rect 9022 2302 9044 2336
rect 9078 2302 9102 2336
rect 9022 2264 9102 2302
rect 9022 2230 9044 2264
rect 9078 2230 9102 2264
rect 9022 2192 9102 2230
rect 9022 2158 9044 2192
rect 9078 2158 9102 2192
rect 9022 2120 9102 2158
rect 9022 2086 9044 2120
rect 9078 2086 9102 2120
rect 9022 2040 9102 2086
rect 9250 2950 9350 3050
rect 9450 2950 9550 3050
rect 9650 2950 9750 3050
rect 9850 2950 9950 3050
rect 10050 2950 10150 3050
rect 10250 2950 10350 3050
rect 10450 2950 10550 3050
rect 10650 2950 10750 3050
rect 10850 2950 10950 3050
rect 9250 2850 10950 2950
rect 9250 2750 9350 2850
rect 9450 2750 9550 2850
rect 9650 2750 9750 2850
rect 9850 2750 9950 2850
rect 10050 2750 10150 2850
rect 10250 2750 10350 2850
rect 10450 2750 10550 2850
rect 10650 2750 10750 2850
rect 10850 2750 10950 2850
rect 9250 2650 10950 2750
rect 9250 2550 9350 2650
rect 9450 2550 9550 2650
rect 9650 2550 9750 2650
rect 9850 2550 9950 2650
rect 10050 2550 10150 2650
rect 10250 2550 10350 2650
rect 10450 2550 10550 2650
rect 10650 2550 10750 2650
rect 10850 2550 10950 2650
rect 9250 2450 10950 2550
rect 9250 2350 9350 2450
rect 9450 2350 9550 2450
rect 9650 2350 9750 2450
rect 9850 2350 9950 2450
rect 10050 2350 10150 2450
rect 10250 2350 10350 2450
rect 10450 2350 10550 2450
rect 10650 2350 10750 2450
rect 10850 2350 10950 2450
rect 9250 2250 10950 2350
rect 9250 2150 9350 2250
rect 9450 2150 9550 2250
rect 9650 2150 9750 2250
rect 9850 2150 9950 2250
rect 10050 2150 10150 2250
rect 10250 2150 10350 2250
rect 10450 2150 10550 2250
rect 10650 2150 10750 2250
rect 10850 2150 10950 2250
rect 9250 2050 10950 2150
rect 9250 1950 9350 2050
rect 9450 1950 9550 2050
rect 9650 1950 9750 2050
rect 9850 1950 9950 2050
rect 10050 1950 10150 2050
rect 10250 1950 10350 2050
rect 10450 1950 10550 2050
rect 10650 1950 10750 2050
rect 10850 1950 10950 2050
rect 11122 2912 11202 2958
rect 11122 2878 11144 2912
rect 11178 2878 11202 2912
rect 11122 2840 11202 2878
rect 11122 2806 11144 2840
rect 11178 2806 11202 2840
rect 11122 2768 11202 2806
rect 11122 2734 11144 2768
rect 11178 2734 11202 2768
rect 11122 2696 11202 2734
rect 11122 2662 11144 2696
rect 11178 2662 11202 2696
rect 11122 2624 11202 2662
rect 11122 2590 11144 2624
rect 11178 2590 11202 2624
rect 11122 2552 11202 2590
rect 11122 2518 11144 2552
rect 11178 2518 11202 2552
rect 11122 2480 11202 2518
rect 11122 2446 11144 2480
rect 11178 2446 11202 2480
rect 11122 2408 11202 2446
rect 11122 2374 11144 2408
rect 11178 2374 11202 2408
rect 11122 2336 11202 2374
rect 11122 2302 11144 2336
rect 11178 2302 11202 2336
rect 11122 2264 11202 2302
rect 11122 2230 11144 2264
rect 11178 2230 11202 2264
rect 11122 2192 11202 2230
rect 11122 2158 11144 2192
rect 11178 2158 11202 2192
rect 11122 2120 11202 2158
rect 11122 2086 11144 2120
rect 11178 2086 11202 2120
rect 11122 2040 11202 2086
rect 13396 2912 13478 2958
rect 13396 2878 13420 2912
rect 13454 2878 13478 2912
rect 13396 2840 13478 2878
rect 13396 2806 13420 2840
rect 13454 2806 13478 2840
rect 13396 2768 13478 2806
rect 13396 2734 13420 2768
rect 13454 2734 13478 2768
rect 13396 2696 13478 2734
rect 13396 2662 13420 2696
rect 13454 2662 13478 2696
rect 13396 2624 13478 2662
rect 13396 2590 13420 2624
rect 13454 2590 13478 2624
rect 13396 2552 13478 2590
rect 13396 2518 13420 2552
rect 13454 2518 13478 2552
rect 13396 2480 13478 2518
rect 13396 2446 13420 2480
rect 13454 2446 13478 2480
rect 13396 2408 13478 2446
rect 13396 2374 13420 2408
rect 13454 2374 13478 2408
rect 13396 2336 13478 2374
rect 13396 2302 13420 2336
rect 13454 2302 13478 2336
rect 13396 2264 13478 2302
rect 13396 2230 13420 2264
rect 13454 2230 13478 2264
rect 13396 2192 13478 2230
rect 13396 2158 13420 2192
rect 13454 2158 13478 2192
rect 13396 2120 13478 2158
rect 13396 2086 13420 2120
rect 13454 2086 13478 2120
rect 13396 2040 13478 2086
rect 13650 2950 13750 3050
rect 13650 2850 13800 2950
rect 13650 2750 13750 2850
rect 13650 2650 13800 2750
rect 13650 2550 13750 2650
rect 13650 2450 13800 2550
rect 13650 2350 13750 2450
rect 13650 2250 13800 2350
rect 13650 2150 13750 2250
rect 13650 2050 13800 2150
rect 13650 1950 13750 2050
rect 0 1850 13800 1950
rect 50 1750 150 1850
rect 250 1750 350 1850
rect 450 1750 550 1850
rect 650 1750 750 1850
rect 850 1750 950 1850
rect 1050 1750 1150 1850
rect 1250 1750 1350 1850
rect 1450 1750 1550 1850
rect 1650 1750 1750 1850
rect 1850 1750 1950 1850
rect 2050 1750 2150 1850
rect 2250 1750 2350 1850
rect 2450 1750 2550 1850
rect 2650 1750 2750 1850
rect 2850 1750 2950 1850
rect 3050 1750 3150 1850
rect 3250 1750 3350 1850
rect 3450 1750 3550 1850
rect 3650 1750 3750 1850
rect 3850 1750 3950 1850
rect 4050 1750 4150 1850
rect 4250 1750 4350 1850
rect 4450 1750 4550 1850
rect 4650 1750 4750 1850
rect 4850 1750 4950 1850
rect 5050 1750 5150 1850
rect 5250 1750 5350 1850
rect 5450 1750 5550 1850
rect 5650 1750 5750 1850
rect 5850 1750 5950 1850
rect 6050 1750 6150 1850
rect 6250 1750 6350 1850
rect 6450 1750 6550 1850
rect 6650 1750 6750 1850
rect 6850 1750 6950 1850
rect 7050 1750 7150 1850
rect 7250 1750 7350 1850
rect 7450 1750 7550 1850
rect 7650 1750 7750 1850
rect 7850 1750 7950 1850
rect 8050 1750 8150 1850
rect 8250 1750 8350 1850
rect 8450 1750 8550 1850
rect 8650 1750 8750 1850
rect 8850 1750 8950 1850
rect 9050 1750 9150 1850
rect 9250 1750 9350 1850
rect 9450 1750 9550 1850
rect 9650 1750 9750 1850
rect 9850 1750 9950 1850
rect 10050 1750 10150 1850
rect 10250 1750 10350 1850
rect 10450 1750 10550 1850
rect 10650 1750 10750 1850
rect 10850 1750 10950 1850
rect 11050 1750 11150 1850
rect 11250 1750 11350 1850
rect 11450 1750 11550 1850
rect 11650 1750 11750 1850
rect 11850 1750 11950 1850
rect 12050 1750 12150 1850
rect 12250 1750 12350 1850
rect 12450 1750 12550 1850
rect 12650 1750 12750 1850
rect 12850 1750 12950 1850
rect 13050 1750 13150 1850
rect 13250 1750 13350 1850
rect 13450 1750 13550 1850
rect 13650 1750 13750 1850
rect 0 1650 13800 1750
rect 50 1550 150 1650
rect 250 1550 350 1650
rect 450 1550 550 1650
rect 650 1550 750 1650
rect 850 1550 950 1650
rect 1050 1550 1150 1650
rect 1250 1550 1350 1650
rect 1450 1550 1550 1650
rect 1650 1550 1750 1650
rect 1850 1550 1950 1650
rect 2050 1550 2150 1650
rect 2250 1550 2350 1650
rect 2450 1550 2550 1650
rect 2650 1550 2750 1650
rect 2850 1550 2950 1650
rect 3050 1550 3150 1650
rect 3250 1550 3350 1650
rect 3450 1550 3550 1650
rect 3650 1550 3750 1650
rect 3850 1550 3950 1650
rect 4050 1550 4150 1650
rect 4250 1550 4350 1650
rect 4450 1550 4550 1650
rect 4650 1550 4750 1650
rect 4850 1550 4950 1650
rect 5050 1550 5150 1650
rect 5250 1550 5350 1650
rect 5450 1550 5550 1650
rect 5650 1550 5750 1650
rect 5850 1550 5950 1650
rect 6050 1550 6150 1650
rect 6250 1550 6350 1650
rect 6450 1550 6550 1650
rect 6650 1550 6750 1650
rect 6850 1550 6950 1650
rect 7050 1550 7150 1650
rect 7250 1550 7350 1650
rect 7450 1550 7550 1650
rect 7650 1550 7750 1650
rect 7850 1550 7950 1650
rect 8050 1550 8150 1650
rect 8250 1550 8350 1650
rect 8450 1550 8550 1650
rect 8650 1550 8750 1650
rect 8850 1550 8950 1650
rect 9050 1550 9150 1650
rect 9250 1550 9350 1650
rect 9450 1550 9550 1650
rect 9650 1550 9750 1650
rect 9850 1550 9950 1650
rect 10050 1550 10150 1650
rect 10250 1550 10350 1650
rect 10450 1550 10550 1650
rect 10650 1550 10750 1650
rect 10850 1550 10950 1650
rect 11050 1550 11150 1650
rect 11250 1550 11350 1650
rect 11450 1550 11550 1650
rect 11650 1550 11750 1650
rect 11850 1550 11950 1650
rect 12050 1550 12150 1650
rect 12250 1550 12350 1650
rect 12450 1550 12550 1650
rect 12650 1550 12750 1650
rect 12850 1550 12950 1650
rect 13050 1550 13150 1650
rect 13250 1550 13350 1650
rect 13450 1550 13550 1650
rect 13650 1550 13750 1650
rect 0 1450 13800 1550
rect 50 1350 150 1450
rect 250 1350 350 1450
rect 450 1350 550 1450
rect 650 1350 750 1450
rect 986 1350 1066 1364
rect 0 1312 1066 1350
rect 0 1278 1008 1312
rect 1042 1278 1066 1312
rect 0 1250 1066 1278
rect 50 1150 150 1250
rect 250 1150 350 1250
rect 450 1150 550 1250
rect 650 1150 750 1250
rect 986 1240 1066 1250
rect 986 1206 1008 1240
rect 1042 1206 1066 1240
rect 986 1168 1066 1206
rect 986 1150 1008 1168
rect 0 1134 1008 1150
rect 1042 1134 1066 1168
rect 0 1096 1066 1134
rect 0 1062 1008 1096
rect 1042 1062 1066 1096
rect 0 1050 1066 1062
rect 50 950 150 1050
rect 250 950 350 1050
rect 450 950 550 1050
rect 650 950 750 1050
rect 986 1024 1066 1050
rect 986 990 1008 1024
rect 1042 990 1066 1024
rect 986 952 1066 990
rect 986 950 1008 952
rect 0 918 1008 950
rect 1042 918 1066 952
rect 0 880 1066 918
rect 0 850 1008 880
rect 50 750 150 850
rect 250 750 350 850
rect 450 750 550 850
rect 650 750 750 850
rect 986 846 1008 850
rect 1042 846 1066 880
rect 986 808 1066 846
rect 986 774 1008 808
rect 1042 774 1066 808
rect 986 750 1066 774
rect 0 736 1066 750
rect 0 702 1008 736
rect 1042 702 1066 736
rect 0 664 1066 702
rect 0 650 1008 664
rect 50 550 150 650
rect 250 550 350 650
rect 450 550 550 650
rect 650 550 750 650
rect 986 630 1008 650
rect 1042 630 1066 664
rect 986 592 1066 630
rect 986 558 1008 592
rect 1042 558 1066 592
rect 986 550 1066 558
rect 0 520 1066 550
rect 0 486 1008 520
rect 1042 486 1066 520
rect 0 450 1066 486
rect 50 350 150 450
rect 250 350 350 450
rect 450 350 550 450
rect 650 350 750 450
rect 986 434 1066 450
rect 6334 1350 6414 1364
rect 6650 1350 6750 1450
rect 6850 1350 6950 1450
rect 7050 1350 7150 1450
rect 7386 1350 7466 1364
rect 6334 1312 7466 1350
rect 6334 1278 6356 1312
rect 6390 1278 7408 1312
rect 7442 1278 7466 1312
rect 6334 1250 7466 1278
rect 6334 1240 6414 1250
rect 6334 1206 6356 1240
rect 6390 1206 6414 1240
rect 6334 1168 6414 1206
rect 6334 1134 6356 1168
rect 6390 1150 6414 1168
rect 6650 1150 6750 1250
rect 6850 1150 6950 1250
rect 7050 1150 7150 1250
rect 7386 1240 7466 1250
rect 7386 1206 7408 1240
rect 7442 1206 7466 1240
rect 7386 1168 7466 1206
rect 7386 1150 7408 1168
rect 6390 1134 7408 1150
rect 7442 1134 7466 1168
rect 6334 1096 7466 1134
rect 6334 1062 6356 1096
rect 6390 1062 7408 1096
rect 7442 1062 7466 1096
rect 6334 1050 7466 1062
rect 6334 1024 6414 1050
rect 6334 990 6356 1024
rect 6390 990 6414 1024
rect 6334 952 6414 990
rect 6334 918 6356 952
rect 6390 950 6414 952
rect 6650 950 6750 1050
rect 6850 950 6950 1050
rect 7050 950 7150 1050
rect 7386 1024 7466 1050
rect 7386 990 7408 1024
rect 7442 990 7466 1024
rect 7386 952 7466 990
rect 7386 950 7408 952
rect 6390 918 7408 950
rect 7442 918 7466 952
rect 6334 880 7466 918
rect 6334 846 6356 880
rect 6390 850 7408 880
rect 6390 846 6414 850
rect 6334 808 6414 846
rect 6334 774 6356 808
rect 6390 774 6414 808
rect 6334 750 6414 774
rect 6650 750 6750 850
rect 6850 750 6950 850
rect 7050 750 7150 850
rect 7386 846 7408 850
rect 7442 846 7466 880
rect 7386 808 7466 846
rect 7386 774 7408 808
rect 7442 774 7466 808
rect 7386 750 7466 774
rect 6334 736 7466 750
rect 6334 702 6356 736
rect 6390 702 7408 736
rect 7442 702 7466 736
rect 6334 664 7466 702
rect 6334 630 6356 664
rect 6390 650 7408 664
rect 6390 630 6414 650
rect 6334 592 6414 630
rect 6334 558 6356 592
rect 6390 558 6414 592
rect 6334 550 6414 558
rect 6650 550 6750 650
rect 6850 550 6950 650
rect 7050 550 7150 650
rect 7386 630 7408 650
rect 7442 630 7466 664
rect 7386 592 7466 630
rect 7386 558 7408 592
rect 7442 558 7466 592
rect 7386 550 7466 558
rect 6334 520 7466 550
rect 6334 486 6356 520
rect 6390 486 7408 520
rect 7442 486 7466 520
rect 6334 450 7466 486
rect 6334 434 6414 450
rect 6650 350 6750 450
rect 6850 350 6950 450
rect 7050 350 7150 450
rect 7386 434 7466 450
rect 12732 1350 12812 1364
rect 13050 1350 13150 1450
rect 13250 1350 13350 1450
rect 13450 1350 13550 1450
rect 13650 1350 13750 1450
rect 12732 1312 13800 1350
rect 12732 1278 12756 1312
rect 12790 1278 13800 1312
rect 12732 1250 13800 1278
rect 12732 1240 12812 1250
rect 12732 1206 12756 1240
rect 12790 1206 12812 1240
rect 12732 1168 12812 1206
rect 12732 1134 12756 1168
rect 12790 1150 12812 1168
rect 13050 1150 13150 1250
rect 13250 1150 13350 1250
rect 13450 1150 13550 1250
rect 13650 1150 13750 1250
rect 12790 1134 13800 1150
rect 12732 1096 13800 1134
rect 12732 1062 12756 1096
rect 12790 1062 13800 1096
rect 12732 1050 13800 1062
rect 12732 1024 12812 1050
rect 12732 990 12756 1024
rect 12790 990 12812 1024
rect 12732 952 12812 990
rect 12732 918 12756 952
rect 12790 950 12812 952
rect 13050 950 13150 1050
rect 13250 950 13350 1050
rect 13450 950 13550 1050
rect 13650 950 13750 1050
rect 12790 918 13800 950
rect 12732 880 13800 918
rect 12732 846 12756 880
rect 12790 850 13800 880
rect 12790 846 12812 850
rect 12732 808 12812 846
rect 12732 774 12756 808
rect 12790 774 12812 808
rect 12732 750 12812 774
rect 13050 750 13150 850
rect 13250 750 13350 850
rect 13450 750 13550 850
rect 13650 750 13750 850
rect 12732 736 13800 750
rect 12732 702 12756 736
rect 12790 702 13800 736
rect 12732 664 13800 702
rect 12732 630 12756 664
rect 12790 650 13800 664
rect 12790 630 12812 650
rect 12732 592 12812 630
rect 12732 558 12756 592
rect 12790 558 12812 592
rect 12732 550 12812 558
rect 13050 550 13150 650
rect 13250 550 13350 650
rect 13450 550 13550 650
rect 13650 550 13750 650
rect 12732 520 13800 550
rect 12732 486 12756 520
rect 12790 486 13800 520
rect 12732 450 13800 486
rect 12732 434 12812 450
rect 13050 350 13150 450
rect 13250 350 13350 450
rect 13450 350 13550 450
rect 13650 350 13750 450
rect 0 250 13800 350
rect 50 150 150 250
rect 250 150 350 250
rect 450 150 550 250
rect 650 150 750 250
rect 850 150 950 250
rect 1050 150 1150 250
rect 1250 150 1350 250
rect 1450 150 1550 250
rect 1650 150 1750 250
rect 1850 150 1950 250
rect 2050 150 2150 250
rect 2250 150 2350 250
rect 2450 150 2550 250
rect 2650 150 2750 250
rect 2850 150 2950 250
rect 3050 150 3150 250
rect 3250 150 3350 250
rect 3450 150 3550 250
rect 3650 150 3750 250
rect 3850 150 3950 250
rect 4050 150 4150 250
rect 4250 150 4350 250
rect 4450 150 4550 250
rect 4650 150 4750 250
rect 4850 150 4950 250
rect 5050 150 5150 250
rect 5250 150 5350 250
rect 5450 150 5550 250
rect 5650 150 5750 250
rect 5850 150 5950 250
rect 6050 150 6150 250
rect 6250 150 6350 250
rect 6450 150 6550 250
rect 6650 150 6750 250
rect 6850 150 6950 250
rect 7050 150 7150 250
rect 7250 150 7350 250
rect 7450 150 7550 250
rect 7650 150 7750 250
rect 7850 150 7950 250
rect 8050 150 8150 250
rect 8250 150 8350 250
rect 8450 150 8550 250
rect 8650 150 8750 250
rect 8850 150 8950 250
rect 9050 150 9150 250
rect 9250 150 9350 250
rect 9450 150 9550 250
rect 9650 150 9750 250
rect 9850 150 9950 250
rect 10050 150 10150 250
rect 10250 150 10350 250
rect 10450 150 10550 250
rect 10650 150 10750 250
rect 10850 150 10950 250
rect 11050 150 11150 250
rect 11250 150 11350 250
rect 11450 150 11550 250
rect 11650 150 11750 250
rect 11850 150 11950 250
rect 12050 150 12150 250
rect 12250 150 12350 250
rect 12450 150 12550 250
rect 12650 150 12750 250
rect 12850 150 12950 250
rect 13050 150 13150 250
rect 13250 150 13350 250
rect 13450 150 13550 250
rect 13650 150 13750 250
rect 0 50 13800 150
rect 50 0 150 50
rect 250 0 350 50
rect 450 0 550 50
rect 650 0 750 50
rect 850 0 950 50
rect 1050 0 1150 50
rect 1250 0 1350 50
rect 1450 0 1550 50
rect 1650 0 1750 50
rect 1850 0 1950 50
rect 2050 0 2150 50
rect 2250 0 2350 50
rect 2450 0 2550 50
rect 2650 0 2750 50
rect 2850 0 2950 50
rect 3050 0 3150 50
rect 3250 0 3350 50
rect 3450 0 3550 50
rect 3650 0 3750 50
rect 3850 0 3950 50
rect 4050 0 4150 50
rect 4250 0 4350 50
rect 4450 0 4550 50
rect 4650 0 4750 50
rect 4850 0 4950 50
rect 5050 0 5150 50
rect 5250 0 5350 50
rect 5450 0 5550 50
rect 5650 0 5750 50
rect 5850 0 5950 50
rect 6050 0 6150 50
rect 6250 0 6350 50
rect 6450 0 6550 50
rect 6650 0 6750 50
rect 6850 0 6950 50
rect 7050 0 7150 50
rect 7250 0 7350 50
rect 7450 0 7550 50
rect 7650 0 7750 50
rect 7850 0 7950 50
rect 8050 0 8150 50
rect 8250 0 8350 50
rect 8450 0 8550 50
rect 8650 0 8750 50
rect 8850 0 8950 50
rect 9050 0 9150 50
rect 9250 0 9350 50
rect 9450 0 9550 50
rect 9650 0 9750 50
rect 9850 0 9950 50
rect 10050 0 10150 50
rect 10250 0 10350 50
rect 10450 0 10550 50
rect 10650 0 10750 50
rect 10850 0 10950 50
rect 11050 0 11150 50
rect 11250 0 11350 50
rect 11450 0 11550 50
rect 11650 0 11750 50
rect 11850 0 11950 50
rect 12050 0 12150 50
rect 12250 0 12350 50
rect 12450 0 12550 50
rect 12650 0 12750 50
rect 12850 0 12950 50
rect 13050 0 13150 50
rect 13250 0 13350 50
rect 13450 0 13550 50
rect 13650 0 13750 50
<< metal2 >>
rect 50 3350 150 3400
rect 250 3350 350 3400
rect 450 3350 550 3400
rect 650 3350 750 3400
rect 850 3350 950 3400
rect 1050 3350 1150 3400
rect 1250 3350 1350 3400
rect 1450 3350 1550 3400
rect 1650 3350 1750 3400
rect 1850 3350 1950 3400
rect 2050 3350 2150 3400
rect 2250 3350 2350 3400
rect 2450 3350 2550 3400
rect 2650 3350 2750 3400
rect 2850 3350 2950 3400
rect 3050 3350 3150 3400
rect 3250 3350 3350 3400
rect 3450 3350 3550 3400
rect 3650 3350 3750 3400
rect 3850 3350 3950 3400
rect 4050 3350 4150 3400
rect 4250 3350 4350 3400
rect 4450 3350 4550 3400
rect 4650 3350 4750 3400
rect 4850 3350 4950 3400
rect 5050 3350 5150 3400
rect 5250 3350 5350 3400
rect 5450 3350 5550 3400
rect 5650 3350 5750 3400
rect 5850 3350 5950 3400
rect 6050 3350 6150 3400
rect 6250 3350 6350 3400
rect 6450 3350 6550 3400
rect 6650 3350 6750 3400
rect 6850 3350 6950 3400
rect 7050 3350 7150 3400
rect 7250 3350 7350 3400
rect 7450 3350 7550 3400
rect 7650 3350 7750 3400
rect 7850 3350 7950 3400
rect 8050 3350 8150 3400
rect 8250 3350 8350 3400
rect 8450 3350 8550 3400
rect 8650 3350 8750 3400
rect 8850 3350 8950 3400
rect 9050 3350 9150 3400
rect 9250 3350 9350 3400
rect 9450 3350 9550 3400
rect 9650 3350 9750 3400
rect 9850 3350 9950 3400
rect 10050 3350 10150 3400
rect 10250 3350 10350 3400
rect 10450 3350 10550 3400
rect 10650 3350 10750 3400
rect 10850 3350 10950 3400
rect 11050 3350 11150 3400
rect 11250 3350 11350 3400
rect 11450 3350 11550 3400
rect 11650 3350 11750 3400
rect 11850 3350 11950 3400
rect 12050 3350 12150 3400
rect 12250 3350 12350 3400
rect 12450 3350 12550 3400
rect 12650 3350 12750 3400
rect 12850 3350 12950 3400
rect 13050 3350 13150 3400
rect 13250 3350 13350 3400
rect 13450 3350 13550 3400
rect 13650 3350 13750 3400
rect 0 3250 13800 3350
rect 50 3150 150 3250
rect 250 3150 350 3250
rect 450 3150 550 3250
rect 650 3150 750 3250
rect 850 3150 950 3250
rect 1050 3150 1150 3250
rect 1250 3150 1350 3250
rect 1450 3150 1550 3250
rect 1650 3150 1750 3250
rect 1850 3150 1950 3250
rect 2050 3150 2150 3250
rect 2250 3150 2350 3250
rect 2450 3150 2550 3250
rect 2650 3150 2750 3250
rect 2850 3150 2950 3250
rect 3050 3150 3150 3250
rect 3250 3150 3350 3250
rect 3450 3150 3550 3250
rect 3650 3150 3750 3250
rect 3850 3150 3950 3250
rect 4050 3150 4150 3250
rect 4250 3150 4350 3250
rect 4450 3150 4550 3250
rect 4650 3150 4750 3250
rect 4850 3150 4950 3250
rect 5050 3150 5150 3250
rect 5250 3150 5350 3250
rect 5450 3150 5550 3250
rect 5650 3150 5750 3250
rect 5850 3150 5950 3250
rect 6050 3150 6150 3250
rect 6250 3150 6350 3250
rect 6450 3150 6550 3250
rect 6650 3150 6750 3250
rect 6850 3150 6950 3250
rect 7050 3150 7150 3250
rect 7250 3150 7350 3250
rect 7450 3150 7550 3250
rect 7650 3150 7750 3250
rect 7850 3150 7950 3250
rect 8050 3150 8150 3250
rect 8250 3150 8350 3250
rect 8450 3150 8550 3250
rect 8650 3150 8750 3250
rect 8850 3150 8950 3250
rect 9050 3150 9150 3250
rect 9250 3150 9350 3250
rect 9450 3150 9550 3250
rect 9650 3150 9750 3250
rect 9850 3150 9950 3250
rect 10050 3150 10150 3250
rect 10250 3150 10350 3250
rect 10450 3150 10550 3250
rect 10650 3150 10750 3250
rect 10850 3150 10950 3250
rect 11050 3150 11150 3250
rect 11250 3150 11350 3250
rect 11450 3150 11550 3250
rect 11650 3150 11750 3250
rect 11850 3150 11950 3250
rect 12050 3150 12150 3250
rect 12250 3150 12350 3250
rect 12450 3150 12550 3250
rect 12650 3150 12750 3250
rect 12850 3150 12950 3250
rect 13050 3150 13150 3250
rect 13250 3150 13350 3250
rect 13450 3150 13550 3250
rect 13650 3150 13750 3250
rect 0 3050 13800 3150
rect 50 2950 150 3050
rect 320 2950 400 2958
rect 0 2850 400 2950
rect 50 2750 150 2850
rect 320 2750 400 2850
rect 0 2650 400 2750
rect 50 2550 150 2650
rect 320 2550 400 2650
rect 0 2450 400 2550
rect 50 2350 150 2450
rect 320 2350 400 2450
rect 0 2250 400 2350
rect 50 2150 150 2250
rect 320 2150 400 2250
rect 0 2050 400 2150
rect 50 1950 150 2050
rect 320 2040 400 2050
rect 2598 2950 2678 2958
rect 2850 2950 2950 3050
rect 3050 2950 3150 3050
rect 3250 2950 3350 3050
rect 3450 2950 3550 3050
rect 3650 2950 3750 3050
rect 3850 2950 3950 3050
rect 4050 2950 4150 3050
rect 4250 2950 4350 3050
rect 4450 2950 4550 3050
rect 4698 2950 4778 2958
rect 2598 2850 4778 2950
rect 2598 2750 2678 2850
rect 2850 2750 2950 2850
rect 3050 2750 3150 2850
rect 3250 2750 3350 2850
rect 3450 2750 3550 2850
rect 3650 2750 3750 2850
rect 3850 2750 3950 2850
rect 4050 2750 4150 2850
rect 4250 2750 4350 2850
rect 4450 2750 4550 2850
rect 4698 2750 4778 2850
rect 2598 2650 4778 2750
rect 2598 2550 2678 2650
rect 2850 2550 2950 2650
rect 3050 2550 3150 2650
rect 3250 2550 3350 2650
rect 3450 2550 3550 2650
rect 3650 2550 3750 2650
rect 3850 2550 3950 2650
rect 4050 2550 4150 2650
rect 4250 2550 4350 2650
rect 4450 2550 4550 2650
rect 4698 2550 4778 2650
rect 2598 2450 4778 2550
rect 2598 2350 2678 2450
rect 2850 2350 2950 2450
rect 3050 2350 3150 2450
rect 3250 2350 3350 2450
rect 3450 2350 3550 2450
rect 3650 2350 3750 2450
rect 3850 2350 3950 2450
rect 4050 2350 4150 2450
rect 4250 2350 4350 2450
rect 4450 2350 4550 2450
rect 4698 2350 4778 2450
rect 2598 2250 4778 2350
rect 2598 2150 2678 2250
rect 2850 2150 2950 2250
rect 3050 2150 3150 2250
rect 3250 2150 3350 2250
rect 3450 2150 3550 2250
rect 3650 2150 3750 2250
rect 3850 2150 3950 2250
rect 4050 2150 4150 2250
rect 4250 2150 4350 2250
rect 4450 2150 4550 2250
rect 4698 2150 4778 2250
rect 2598 2050 4778 2150
rect 2598 2040 2678 2050
rect 2850 1950 2950 2050
rect 3050 1950 3150 2050
rect 3250 1950 3350 2050
rect 3450 1950 3550 2050
rect 3650 1950 3750 2050
rect 3850 1950 3950 2050
rect 4050 1950 4150 2050
rect 4250 1950 4350 2050
rect 4450 1950 4550 2050
rect 4698 2040 4778 2050
rect 9022 2950 9102 2958
rect 9250 2950 9350 3050
rect 9450 2950 9550 3050
rect 9650 2950 9750 3050
rect 9850 2950 9950 3050
rect 10050 2950 10150 3050
rect 10250 2950 10350 3050
rect 10450 2950 10550 3050
rect 10650 2950 10750 3050
rect 10850 2950 10950 3050
rect 11122 2950 11202 2958
rect 9022 2850 11202 2950
rect 9022 2750 9102 2850
rect 9250 2750 9350 2850
rect 9450 2750 9550 2850
rect 9650 2750 9750 2850
rect 9850 2750 9950 2850
rect 10050 2750 10150 2850
rect 10250 2750 10350 2850
rect 10450 2750 10550 2850
rect 10650 2750 10750 2850
rect 10850 2750 10950 2850
rect 11122 2750 11202 2850
rect 9022 2650 11202 2750
rect 9022 2550 9102 2650
rect 9250 2550 9350 2650
rect 9450 2550 9550 2650
rect 9650 2550 9750 2650
rect 9850 2550 9950 2650
rect 10050 2550 10150 2650
rect 10250 2550 10350 2650
rect 10450 2550 10550 2650
rect 10650 2550 10750 2650
rect 10850 2550 10950 2650
rect 11122 2550 11202 2650
rect 9022 2450 11202 2550
rect 9022 2350 9102 2450
rect 9250 2350 9350 2450
rect 9450 2350 9550 2450
rect 9650 2350 9750 2450
rect 9850 2350 9950 2450
rect 10050 2350 10150 2450
rect 10250 2350 10350 2450
rect 10450 2350 10550 2450
rect 10650 2350 10750 2450
rect 10850 2350 10950 2450
rect 11122 2350 11202 2450
rect 9022 2250 11202 2350
rect 9022 2150 9102 2250
rect 9250 2150 9350 2250
rect 9450 2150 9550 2250
rect 9650 2150 9750 2250
rect 9850 2150 9950 2250
rect 10050 2150 10150 2250
rect 10250 2150 10350 2250
rect 10450 2150 10550 2250
rect 10650 2150 10750 2250
rect 10850 2150 10950 2250
rect 11122 2150 11202 2250
rect 9022 2050 11202 2150
rect 9022 2040 9102 2050
rect 9250 1950 9350 2050
rect 9450 1950 9550 2050
rect 9650 1950 9750 2050
rect 9850 1950 9950 2050
rect 10050 1950 10150 2050
rect 10250 1950 10350 2050
rect 10450 1950 10550 2050
rect 10650 1950 10750 2050
rect 10850 1950 10950 2050
rect 11122 2040 11202 2050
rect 13396 2950 13478 2958
rect 13650 2950 13750 3050
rect 13396 2850 13800 2950
rect 13396 2750 13478 2850
rect 13650 2750 13750 2850
rect 13396 2650 13800 2750
rect 13396 2550 13478 2650
rect 13650 2550 13750 2650
rect 13396 2450 13800 2550
rect 13396 2350 13478 2450
rect 13650 2350 13750 2450
rect 13396 2250 13800 2350
rect 13396 2150 13478 2250
rect 13650 2150 13750 2250
rect 13396 2050 13800 2150
rect 13396 2040 13478 2050
rect 13650 1950 13750 2050
rect 0 1850 13800 1950
rect 50 1750 150 1850
rect 250 1750 350 1850
rect 450 1750 550 1850
rect 650 1750 750 1850
rect 850 1750 950 1850
rect 1050 1750 1150 1850
rect 1250 1750 1350 1850
rect 1450 1750 1550 1850
rect 1650 1750 1750 1850
rect 1850 1750 1950 1850
rect 2050 1750 2150 1850
rect 2250 1750 2350 1850
rect 2450 1750 2550 1850
rect 2650 1750 2750 1850
rect 2850 1750 2950 1850
rect 3050 1750 3150 1850
rect 3250 1750 3350 1850
rect 3450 1750 3550 1850
rect 3650 1750 3750 1850
rect 3850 1750 3950 1850
rect 4050 1750 4150 1850
rect 4250 1750 4350 1850
rect 4450 1750 4550 1850
rect 4650 1750 4750 1850
rect 4850 1750 4950 1850
rect 5050 1750 5150 1850
rect 5250 1750 5350 1850
rect 5450 1750 5550 1850
rect 5650 1750 5750 1850
rect 5850 1750 5950 1850
rect 6050 1750 6150 1850
rect 6250 1750 6350 1850
rect 6450 1750 6550 1850
rect 6650 1750 6750 1850
rect 6850 1750 6950 1850
rect 7050 1750 7150 1850
rect 7250 1750 7350 1850
rect 7450 1750 7550 1850
rect 7650 1750 7750 1850
rect 7850 1750 7950 1850
rect 8050 1750 8150 1850
rect 8250 1750 8350 1850
rect 8450 1750 8550 1850
rect 8650 1750 8750 1850
rect 8850 1750 8950 1850
rect 9050 1750 9150 1850
rect 9250 1750 9350 1850
rect 9450 1750 9550 1850
rect 9650 1750 9750 1850
rect 9850 1750 9950 1850
rect 10050 1750 10150 1850
rect 10250 1750 10350 1850
rect 10450 1750 10550 1850
rect 10650 1750 10750 1850
rect 10850 1750 10950 1850
rect 11050 1750 11150 1850
rect 11250 1750 11350 1850
rect 11450 1750 11550 1850
rect 11650 1750 11750 1850
rect 11850 1750 11950 1850
rect 12050 1750 12150 1850
rect 12250 1750 12350 1850
rect 12450 1750 12550 1850
rect 12650 1750 12750 1850
rect 12850 1750 12950 1850
rect 13050 1750 13150 1850
rect 13250 1750 13350 1850
rect 13450 1750 13550 1850
rect 13650 1750 13750 1850
rect 0 1650 13800 1750
rect 50 1550 150 1650
rect 250 1550 350 1650
rect 450 1550 550 1650
rect 650 1550 750 1650
rect 850 1550 950 1650
rect 1050 1550 1150 1650
rect 1250 1550 1350 1650
rect 1450 1550 1550 1650
rect 1650 1550 1750 1650
rect 1850 1550 1950 1650
rect 2050 1550 2150 1650
rect 2250 1550 2350 1650
rect 2450 1550 2550 1650
rect 2650 1550 2750 1650
rect 2850 1550 2950 1650
rect 3050 1550 3150 1650
rect 3250 1550 3350 1650
rect 3450 1550 3550 1650
rect 3650 1550 3750 1650
rect 3850 1550 3950 1650
rect 4050 1550 4150 1650
rect 4250 1550 4350 1650
rect 4450 1550 4550 1650
rect 4650 1550 4750 1650
rect 4850 1550 4950 1650
rect 5050 1550 5150 1650
rect 5250 1550 5350 1650
rect 5450 1550 5550 1650
rect 5650 1550 5750 1650
rect 5850 1550 5950 1650
rect 6050 1550 6150 1650
rect 6250 1550 6350 1650
rect 6450 1550 6550 1650
rect 6650 1550 6750 1650
rect 6850 1550 6950 1650
rect 7050 1550 7150 1650
rect 7250 1550 7350 1650
rect 7450 1550 7550 1650
rect 7650 1550 7750 1650
rect 7850 1550 7950 1650
rect 8050 1550 8150 1650
rect 8250 1550 8350 1650
rect 8450 1550 8550 1650
rect 8650 1550 8750 1650
rect 8850 1550 8950 1650
rect 9050 1550 9150 1650
rect 9250 1550 9350 1650
rect 9450 1550 9550 1650
rect 9650 1550 9750 1650
rect 9850 1550 9950 1650
rect 10050 1550 10150 1650
rect 10250 1550 10350 1650
rect 10450 1550 10550 1650
rect 10650 1550 10750 1650
rect 10850 1550 10950 1650
rect 11050 1550 11150 1650
rect 11250 1550 11350 1650
rect 11450 1550 11550 1650
rect 11650 1550 11750 1650
rect 11850 1550 11950 1650
rect 12050 1550 12150 1650
rect 12250 1550 12350 1650
rect 12450 1550 12550 1650
rect 12650 1550 12750 1650
rect 12850 1550 12950 1650
rect 13050 1550 13150 1650
rect 13250 1550 13350 1650
rect 13450 1550 13550 1650
rect 13650 1550 13750 1650
rect 0 1450 13800 1550
rect 50 1350 150 1450
rect 250 1350 350 1450
rect 450 1350 550 1450
rect 650 1350 750 1450
rect 0 1250 750 1350
rect 50 1150 150 1250
rect 250 1150 350 1250
rect 450 1150 550 1250
rect 650 1150 750 1250
rect 0 1050 750 1150
rect 50 950 150 1050
rect 250 950 350 1050
rect 450 950 550 1050
rect 650 950 750 1050
rect 0 850 750 950
rect 50 750 150 850
rect 250 750 350 850
rect 450 750 550 850
rect 650 750 750 850
rect 0 650 750 750
rect 50 550 150 650
rect 250 550 350 650
rect 450 550 550 650
rect 650 550 750 650
rect 0 450 750 550
rect 50 350 150 450
rect 250 350 350 450
rect 450 350 550 450
rect 650 350 750 450
rect 6650 1350 6750 1450
rect 6850 1350 6950 1450
rect 7050 1350 7150 1450
rect 6650 1250 7150 1350
rect 6650 1150 6750 1250
rect 6850 1150 6950 1250
rect 7050 1150 7150 1250
rect 6650 1050 7150 1150
rect 6650 950 6750 1050
rect 6850 950 6950 1050
rect 7050 950 7150 1050
rect 6650 850 7150 950
rect 6650 750 6750 850
rect 6850 750 6950 850
rect 7050 750 7150 850
rect 6650 650 7150 750
rect 6650 550 6750 650
rect 6850 550 6950 650
rect 7050 550 7150 650
rect 6650 450 7150 550
rect 6650 350 6750 450
rect 6850 350 6950 450
rect 7050 350 7150 450
rect 13050 1350 13150 1450
rect 13250 1350 13350 1450
rect 13450 1350 13550 1450
rect 13650 1350 13750 1450
rect 13050 1250 13800 1350
rect 13050 1150 13150 1250
rect 13250 1150 13350 1250
rect 13450 1150 13550 1250
rect 13650 1150 13750 1250
rect 13050 1050 13800 1150
rect 13050 950 13150 1050
rect 13250 950 13350 1050
rect 13450 950 13550 1050
rect 13650 950 13750 1050
rect 13050 850 13800 950
rect 13050 750 13150 850
rect 13250 750 13350 850
rect 13450 750 13550 850
rect 13650 750 13750 850
rect 13050 650 13800 750
rect 13050 550 13150 650
rect 13250 550 13350 650
rect 13450 550 13550 650
rect 13650 550 13750 650
rect 13050 450 13800 550
rect 13050 350 13150 450
rect 13250 350 13350 450
rect 13450 350 13550 450
rect 13650 350 13750 450
rect 0 250 13800 350
rect 50 150 150 250
rect 250 150 350 250
rect 450 150 550 250
rect 650 150 750 250
rect 850 150 950 250
rect 1050 150 1150 250
rect 1250 150 1350 250
rect 1450 150 1550 250
rect 1650 150 1750 250
rect 1850 150 1950 250
rect 2050 150 2150 250
rect 2250 150 2350 250
rect 2450 150 2550 250
rect 2650 150 2750 250
rect 2850 150 2950 250
rect 3050 150 3150 250
rect 3250 150 3350 250
rect 3450 150 3550 250
rect 3650 150 3750 250
rect 3850 150 3950 250
rect 4050 150 4150 250
rect 4250 150 4350 250
rect 4450 150 4550 250
rect 4650 150 4750 250
rect 4850 150 4950 250
rect 5050 150 5150 250
rect 5250 150 5350 250
rect 5450 150 5550 250
rect 5650 150 5750 250
rect 5850 150 5950 250
rect 6050 150 6150 250
rect 6250 150 6350 250
rect 6450 150 6550 250
rect 6650 150 6750 250
rect 6850 150 6950 250
rect 7050 150 7150 250
rect 7250 150 7350 250
rect 7450 150 7550 250
rect 7650 150 7750 250
rect 7850 150 7950 250
rect 8050 150 8150 250
rect 8250 150 8350 250
rect 8450 150 8550 250
rect 8650 150 8750 250
rect 8850 150 8950 250
rect 9050 150 9150 250
rect 9250 150 9350 250
rect 9450 150 9550 250
rect 9650 150 9750 250
rect 9850 150 9950 250
rect 10050 150 10150 250
rect 10250 150 10350 250
rect 10450 150 10550 250
rect 10650 150 10750 250
rect 10850 150 10950 250
rect 11050 150 11150 250
rect 11250 150 11350 250
rect 11450 150 11550 250
rect 11650 150 11750 250
rect 11850 150 11950 250
rect 12050 150 12150 250
rect 12250 150 12350 250
rect 12450 150 12550 250
rect 12650 150 12750 250
rect 12850 150 12950 250
rect 13050 150 13150 250
rect 13250 150 13350 250
rect 13450 150 13550 250
rect 13650 150 13750 250
rect 0 50 13800 150
rect 50 0 150 50
rect 250 0 350 50
rect 450 0 550 50
rect 650 0 750 50
rect 850 0 950 50
rect 1050 0 1150 50
rect 1250 0 1350 50
rect 1450 0 1550 50
rect 1650 0 1750 50
rect 1850 0 1950 50
rect 2050 0 2150 50
rect 2250 0 2350 50
rect 2450 0 2550 50
rect 2650 0 2750 50
rect 2850 0 2950 50
rect 3050 0 3150 50
rect 3250 0 3350 50
rect 3450 0 3550 50
rect 3650 0 3750 50
rect 3850 0 3950 50
rect 4050 0 4150 50
rect 4250 0 4350 50
rect 4450 0 4550 50
rect 4650 0 4750 50
rect 4850 0 4950 50
rect 5050 0 5150 50
rect 5250 0 5350 50
rect 5450 0 5550 50
rect 5650 0 5750 50
rect 5850 0 5950 50
rect 6050 0 6150 50
rect 6250 0 6350 50
rect 6450 0 6550 50
rect 6650 0 6750 50
rect 6850 0 6950 50
rect 7050 0 7150 50
rect 7250 0 7350 50
rect 7450 0 7550 50
rect 7650 0 7750 50
rect 7850 0 7950 50
rect 8050 0 8150 50
rect 8250 0 8350 50
rect 8450 0 8550 50
rect 8650 0 8750 50
rect 8850 0 8950 50
rect 9050 0 9150 50
rect 9250 0 9350 50
rect 9450 0 9550 50
rect 9650 0 9750 50
rect 9850 0 9950 50
rect 10050 0 10150 50
rect 10250 0 10350 50
rect 10450 0 10550 50
rect 10650 0 10750 50
rect 10850 0 10950 50
rect 11050 0 11150 50
rect 11250 0 11350 50
rect 11450 0 11550 50
rect 11650 0 11750 50
rect 11850 0 11950 50
rect 12050 0 12150 50
rect 12250 0 12350 50
rect 12450 0 12550 50
rect 12650 0 12750 50
rect 12850 0 12950 50
rect 13050 0 13150 50
rect 13250 0 13350 50
rect 13450 0 13550 50
rect 13650 0 13750 50
<< metal3 >>
rect 1850 2450 1950 2550
rect 2250 2540 2350 2550
rect 4850 2540 4950 2550
rect 2250 2460 4950 2540
rect 2250 2450 2350 2460
rect 4850 2450 4950 2460
rect 8850 2540 8950 2550
rect 11450 2540 11550 2550
rect 8850 2460 11550 2540
rect 8850 2450 8950 2460
rect 11450 2450 11550 2460
rect 11850 2450 11950 2550
rect 2250 2050 2350 2150
rect 11450 2050 11550 2150
rect 1850 1250 1950 1350
rect 3650 1250 3750 1350
rect 6050 1340 6150 1350
rect 7650 1340 7750 1350
rect 6050 1260 7750 1340
rect 6050 1250 6150 1260
rect 7650 1250 7750 1260
rect 3650 850 3750 950
rect 11850 850 11950 950
<< metal4 >>
rect 1860 1260 1940 2540
rect 2260 2060 2340 2540
rect 11460 2060 11540 2540
rect 3660 860 3740 1340
rect 11860 860 11940 2540
use via_M1_M2_1_a  NoName_294 ~/A2G/MAGIC/magic_layout/skywater130_microtemplates_dense
timestamp 1647525606
transform 1 0 360 0 1 2500
box -32 -32 32 32
use via_M1_M2_1_b  NoName_295 ~/A2G/MAGIC/magic_layout/skywater130_microtemplates_dense
timestamp 1647525606
transform 1 0 360 0 1 2628
box -32 -32 32 32
use via_M1_M2_1_c  NoName_296 ~/A2G/MAGIC/magic_layout/skywater130_microtemplates_dense
timestamp 1647525606
transform 1 0 360 0 1 2372
box -32 -32 32 32
use via_M1_M2_1_d  NoName_297 ~/A2G/MAGIC/magic_layout/skywater130_microtemplates_dense
timestamp 1647525606
transform 1 0 360 0 1 2756
box -32 -32 32 32
use via_M1_M2_1_e  NoName_298 ~/A2G/MAGIC/magic_layout/skywater130_microtemplates_dense
timestamp 1647525606
transform 1 0 360 0 1 2244
box -32 -32 32 32
use via_M1_M2_1_f  NoName_299 ~/A2G/MAGIC/magic_layout/skywater130_microtemplates_dense
timestamp 1647525606
transform 1 0 360 0 1 2884
box -32 -32 32 32
use via_M1_M2_1_g  NoName_300 ~/A2G/MAGIC/magic_layout/skywater130_microtemplates_dense
timestamp 1647525606
transform 1 0 360 0 1 2116
box -32 -32 32 32
use via_M1_M2_1_h  NoName_301 ~/A2G/MAGIC/magic_layout/skywater130_microtemplates_dense
timestamp 1647525606
transform 1 0 2638 0 1 2500
box -32 -32 32 32
use via_M1_M2_1_i  NoName_302 ~/A2G/MAGIC/magic_layout/skywater130_microtemplates_dense
timestamp 1647525606
transform 1 0 2638 0 1 2628
box -32 -32 32 32
use via_M1_M2_1_j  NoName_303 ~/A2G/MAGIC/magic_layout/skywater130_microtemplates_dense
timestamp 1647525606
transform 1 0 2638 0 1 2372
box -32 -32 32 32
use via_M1_M2_1_k  NoName_304 ~/A2G/MAGIC/magic_layout/skywater130_microtemplates_dense
timestamp 1647525606
transform 1 0 2638 0 1 2756
box -32 -32 32 32
use via_M1_M2_1_l  NoName_305 ~/A2G/MAGIC/magic_layout/skywater130_microtemplates_dense
timestamp 1647525606
transform 1 0 2638 0 1 2244
box -32 -32 32 32
use via_M1_M2_1_m  NoName_306 ~/A2G/MAGIC/magic_layout/skywater130_microtemplates_dense
timestamp 1647525606
transform 1 0 2638 0 1 2884
box -32 -32 32 32
use via_M1_M2_1_n  NoName_307 ~/A2G/MAGIC/magic_layout/skywater130_microtemplates_dense
timestamp 1647525606
transform 1 0 2638 0 1 2116
box -32 -32 32 32
use via_M1_M2_1_o  NoName_308 ~/A2G/MAGIC/magic_layout/skywater130_microtemplates_dense
timestamp 1647525606
transform 1 0 11162 0 1 2500
box -32 -32 32 32
use via_M1_M2_1_p  NoName_309 ~/A2G/MAGIC/magic_layout/skywater130_microtemplates_dense
timestamp 1647525606
transform 1 0 11162 0 1 2628
box -32 -32 32 32
use via_M1_M2_1_q  NoName_310 ~/A2G/MAGIC/magic_layout/skywater130_microtemplates_dense
timestamp 1647525606
transform 1 0 11162 0 1 2372
box -32 -32 32 32
use via_M1_M2_1_r  NoName_311 ~/A2G/MAGIC/magic_layout/skywater130_microtemplates_dense
timestamp 1647525606
transform 1 0 11162 0 1 2756
box -32 -32 32 32
use via_M1_M2_1_s  NoName_312 ~/A2G/MAGIC/magic_layout/skywater130_microtemplates_dense
timestamp 1647525606
transform 1 0 11162 0 1 2244
box -32 -32 32 32
use via_M1_M2_1_t  NoName_313 ~/A2G/MAGIC/magic_layout/skywater130_microtemplates_dense
timestamp 1647525606
transform 1 0 11162 0 1 2884
box -32 -32 32 32
use via_M1_M2_1_u  NoName_314 ~/A2G/MAGIC/magic_layout/skywater130_microtemplates_dense
timestamp 1647525606
transform 1 0 11162 0 1 2116
box -32 -32 32 32
use via_M1_M2_1_v  NoName_315 ~/A2G/MAGIC/magic_layout/skywater130_microtemplates_dense
timestamp 1647525606
transform 1 0 13438 0 1 2500
box -32 -32 32 32
use via_M1_M2_1_w  NoName_316 ~/A2G/MAGIC/magic_layout/skywater130_microtemplates_dense
timestamp 1647525606
transform 1 0 13438 0 1 2628
box -32 -32 32 32
use via_M1_M2_1_x  NoName_317 ~/A2G/MAGIC/magic_layout/skywater130_microtemplates_dense
timestamp 1647525606
transform 1 0 13438 0 1 2372
box -32 -32 32 32
use via_M1_M2_1_y  NoName_318 ~/A2G/MAGIC/magic_layout/skywater130_microtemplates_dense
timestamp 1647525606
transform 1 0 13438 0 1 2756
box -32 -32 32 32
use via_M1_M2_1_z  NoName_319 ~/A2G/MAGIC/magic_layout/skywater130_microtemplates_dense
timestamp 1647525606
transform 1 0 13438 0 1 2244
box -32 -32 32 32
use via_M1_M2_1_{  NoName_320 ~/A2G/MAGIC/magic_layout/skywater130_microtemplates_dense
timestamp 1647525606
transform 1 0 13438 0 1 2884
box -32 -32 32 32
use via_M1_M2_1_|  NoName_321 ~/A2G/MAGIC/magic_layout/skywater130_microtemplates_dense
timestamp 1647525606
transform 1 0 13438 0 1 2116
box -32 -32 32 32
use via_M1_M2_1_}  NoName_322 ~/A2G/MAGIC/magic_layout/skywater130_microtemplates_dense
timestamp 1647525606
transform 1 0 4738 0 1 2500
box -32 -32 32 32
use via_M1_M2_1_~  NoName_323 ~/A2G/MAGIC/magic_layout/skywater130_microtemplates_dense
timestamp 1647525606
transform 1 0 4738 0 1 2628
box -32 -32 32 32
use via_M1_M2_1_  NoName_324 ~/A2G/MAGIC/magic_layout/skywater130_microtemplates_dense
timestamp 1647525606
transform 1 0 4738 0 1 2372
box -32 -32 32 32
use via_M1_M2_1_�  NoName_325 ~/A2G/MAGIC/magic_layout/skywater130_microtemplates_dense
timestamp 1647525606
transform 1 0 4738 0 1 2756
box -32 -32 32 32
use via_M1_M2_1_�  NoName_326 ~/A2G/MAGIC/magic_layout/skywater130_microtemplates_dense
timestamp 1647525606
transform 1 0 4738 0 1 2244
box -32 -32 32 32
use via_M1_M2_1_�  NoName_327 ~/A2G/MAGIC/magic_layout/skywater130_microtemplates_dense
timestamp 1647525606
transform 1 0 4738 0 1 2884
box -32 -32 32 32
use via_M1_M2_1_�  NoName_328 ~/A2G/MAGIC/magic_layout/skywater130_microtemplates_dense
timestamp 1647525606
transform 1 0 4738 0 1 2116
box -32 -32 32 32
use via_M1_M2_1_�  NoName_329 ~/A2G/MAGIC/magic_layout/skywater130_microtemplates_dense
timestamp 1647525606
transform 1 0 9062 0 1 2500
box -32 -32 32 32
use via_M1_M2_1_�  NoName_330 ~/A2G/MAGIC/magic_layout/skywater130_microtemplates_dense
timestamp 1647525606
transform 1 0 9062 0 1 2628
box -32 -32 32 32
use via_M1_M2_1_�  NoName_331 ~/A2G/MAGIC/magic_layout/skywater130_microtemplates_dense
timestamp 1647525606
transform 1 0 9062 0 1 2372
box -32 -32 32 32
use via_M1_M2_1_�  NoName_332 ~/A2G/MAGIC/magic_layout/skywater130_microtemplates_dense
timestamp 1647525606
transform 1 0 9062 0 1 2756
box -32 -32 32 32
use via_M1_M2_1_�  NoName_333 ~/A2G/MAGIC/magic_layout/skywater130_microtemplates_dense
timestamp 1647525606
transform 1 0 9062 0 1 2244
box -32 -32 32 32
use via_M1_M2_1_�  NoName_334 ~/A2G/MAGIC/magic_layout/skywater130_microtemplates_dense
timestamp 1647525606
transform 1 0 9062 0 1 2884
box -32 -32 32 32
use via_M1_M2_1_�  NoName_335 ~/A2G/MAGIC/magic_layout/skywater130_microtemplates_dense
timestamp 1647525606
transform 1 0 9062 0 1 2116
box -32 -32 32 32
use via_M2_M3_0  NoName_336 ~/A2G/MAGIC/magic_layout/skywater130_microtemplates_dense
timestamp 1647525786
transform 1 0 3700 0 1 900
box -38 -38 38 38
use via_M2_M3_0  NoName_337
timestamp 1647525786
transform 1 0 3700 0 1 1300
box -38 -38 38 38
use via_M3_M4_0  NoName_339 ~/A2G/MAGIC/magic_layout/skywater130_microtemplates_dense
timestamp 1647526059
transform 1 0 3700 0 1 900
box -38 -38 38 38
use via_M3_M4_0  NoName_340
timestamp 1647526059
transform 1 0 3700 0 1 1300
box -38 -38 38 38
use via_M2_M3_0  NoName_342
timestamp 1647525786
transform 1 0 1900 0 1 2500
box -38 -38 38 38
use via_M2_M3_0  NoName_343
timestamp 1647525786
transform 1 0 1900 0 1 1300
box -38 -38 38 38
use via_M3_M4_0  NoName_345
timestamp 1647526059
transform 1 0 1900 0 1 2500
box -38 -38 38 38
use via_M3_M4_0  NoName_346
timestamp 1647526059
transform 1 0 1900 0 1 1300
box -38 -38 38 38
use via_M2_M3_0  NoName_348
timestamp 1647525786
transform 1 0 6100 0 1 1300
box -38 -38 38 38
use via_M2_M3_0  NoName_349
timestamp 1647525786
transform 1 0 7700 0 1 1300
box -38 -38 38 38
use via_M2_M3_0  NoName_352
timestamp 1647525786
transform 1 0 2300 0 1 2100
box -38 -38 38 38
use via_M2_M3_0  NoName_353
timestamp 1647525786
transform 1 0 4900 0 1 2500
box -38 -38 38 38
use via_M3_M4_0  NoName_355
timestamp 1647526059
transform 1 0 2300 0 1 2100
box -38 -38 38 38
use via_M3_M4_0  NoName_356
timestamp 1647526059
transform 1 0 2300 0 1 2500
box -38 -38 38 38
use via_M2_M3_0  NoName_358
timestamp 1647525786
transform 1 0 11500 0 1 2100
box -38 -38 38 38
use via_M2_M3_0  NoName_359
timestamp 1647525786
transform 1 0 8900 0 1 2500
box -38 -38 38 38
use via_M3_M4_0  NoName_361
timestamp 1647526059
transform 1 0 11500 0 1 2100
box -38 -38 38 38
use via_M3_M4_0  NoName_362
timestamp 1647526059
transform 1 0 11500 0 1 2500
box -38 -38 38 38
use via_M2_M3_0  NoName_364
timestamp 1647525786
transform 1 0 11900 0 1 2500
box -38 -38 38 38
use via_M2_M3_0  NoName_365
timestamp 1647525786
transform 1 0 11900 0 1 900
box -38 -38 38 38
use via_M3_M4_0  NoName_367
timestamp 1647526059
transform 1 0 11900 0 1 2500
box -38 -38 38 38
use via_M3_M4_0  NoName_368
timestamp 1647526059
transform 1 0 11900 0 1 900
box -38 -38 38 38
use XM1  XM1 ~/A2G/MAGIC/magic_layout/pcell
timestamp 1679394721
transform 1 0 1500 0 1 2500
box -1191 -529 1191 529
use XM2  XM2 ~/A2G/MAGIC/magic_layout/pcell
timestamp 1679394722
transform 1 0 3700 0 1 900
box -2727 -534 2727 534
use XM3  XM3 ~/A2G/MAGIC/magic_layout/pcell
timestamp 1679394722
transform 1 0 12300 0 1 2500
box -1191 -529 1191 529
use XM4  XM4 ~/A2G/MAGIC/magic_layout/pcell
timestamp 1679394723
transform 1 0 10100 0 1 900
box -2727 -534 2727 534
use XM5  XM5 ~/A2G/MAGIC/magic_layout/pcell
timestamp 1679394724
transform 1 0 6900 0 1 2500
box -2215 -529 2215 529
<< labels >>
flabel metal3 3700 900 3700 900 0 FreeSans 1600 0 0 0 XM2_D
flabel metal4 3700 1300 3700 1300 0 FreeSans 1600 0 0 0 XM2_G
flabel metal3 1900 2500 1900 2500 0 FreeSans 1600 0 0 0 XM1_D
flabel metal4 1900 1300 1900 1300 0 FreeSans 1600 0 0 0 XM2_G
flabel metal3 6100 1300 6100 1300 0 FreeSans 1600 0 0 0 XM2_G
flabel metal3 7700 1300 7700 1300 0 FreeSans 1600 0 0 0 XM4_G
flabel metal3 2300 2100 2300 2100 0 FreeSans 1600 0 0 0 XM1_S
flabel metal3 4900 2500 4900 2500 0 FreeSans 1600 0 0 0 XM5_D
flabel metal3 11500 2100 11500 2100 0 FreeSans 1600 0 0 0 XM3_S
flabel metal3 8900 2500 8900 2500 0 FreeSans 1600 0 0 0 XM5_D
flabel metal3 11900 2500 11900 2500 0 FreeSans 1600 0 0 0 XM3_D
flabel metal4 11900 900 11900 900 0 FreeSans 1600 0 0 0 XM4_D
flabel metal3 1500 2900 1500 2900 0 FreeSans 1600 0 0 0 ia
flabel metal3 6900 2100 6900 2100 0 FreeSans 1600 0 0 0 vss
flabel metal3 3700 500 3700 500 0 FreeSans 1600 0 0 0 vdd
flabel metal3 10100 500 10100 500 0 FreeSans 1600 0 0 0 vdd
flabel metal3 12300 2900 12300 2900 0 FreeSans 1600 0 0 0 ib
flabel metal3 6900 2900 6900 2900 0 FreeSans 1600 0 0 0 icmbias
<< end >>
