magic
tech sky130A
magscale 1 2
timestamp 1686266346
<< checkpaint >>
rect -2135 -1799 2135 1799
<< pwell >>
rect -875 -539 875 539
<< nmos >>
rect -679 -391 -619 329
rect -561 -391 -501 329
rect -443 -391 -383 329
rect -325 -391 -265 329
rect -207 -391 -147 329
rect -89 -391 -29 329
rect 29 -391 89 329
rect 147 -391 207 329
rect 265 -391 325 329
rect 383 -391 443 329
rect 501 -391 561 329
rect 619 -391 679 329
<< ndiff >>
rect -737 317 -679 329
rect -737 -379 -725 317
rect -691 -379 -679 317
rect -737 -391 -679 -379
rect -619 317 -561 329
rect -619 -379 -607 317
rect -573 -379 -561 317
rect -619 -391 -561 -379
rect -501 317 -443 329
rect -501 -379 -489 317
rect -455 -379 -443 317
rect -501 -391 -443 -379
rect -383 317 -325 329
rect -383 -379 -371 317
rect -337 -379 -325 317
rect -383 -391 -325 -379
rect -265 317 -207 329
rect -265 -379 -253 317
rect -219 -379 -207 317
rect -265 -391 -207 -379
rect -147 317 -89 329
rect -147 -379 -135 317
rect -101 -379 -89 317
rect -147 -391 -89 -379
rect -29 317 29 329
rect -29 -379 -17 317
rect 17 -379 29 317
rect -29 -391 29 -379
rect 89 317 147 329
rect 89 -379 101 317
rect 135 -379 147 317
rect 89 -391 147 -379
rect 207 317 265 329
rect 207 -379 219 317
rect 253 -379 265 317
rect 207 -391 265 -379
rect 325 317 383 329
rect 325 -379 337 317
rect 371 -379 383 317
rect 325 -391 383 -379
rect 443 317 501 329
rect 443 -379 455 317
rect 489 -379 501 317
rect 443 -391 501 -379
rect 561 317 619 329
rect 561 -379 573 317
rect 607 -379 619 317
rect 561 -391 619 -379
rect 679 317 737 329
rect 679 -379 691 317
rect 725 -379 737 317
rect 679 -391 737 -379
<< ndiffc >>
rect -725 -379 -691 317
rect -607 -379 -573 317
rect -489 -379 -455 317
rect -371 -379 -337 317
rect -253 -379 -219 317
rect -135 -379 -101 317
rect -17 -379 17 317
rect 101 -379 135 317
rect 219 -379 253 317
rect 337 -379 371 317
rect 455 -379 489 317
rect 573 -379 607 317
rect 691 -379 725 317
<< psubdiff >>
rect -839 469 -743 503
rect 743 469 839 503
rect -839 407 -805 469
rect 805 407 839 469
rect -839 -469 -805 -407
rect 805 -469 839 -407
rect -839 -503 -743 -469
rect 743 -503 839 -469
<< psubdiffcont >>
rect -743 469 743 503
rect -839 -407 -805 407
rect 805 -407 839 407
rect -743 -503 743 -469
<< poly >>
rect -682 401 -616 417
rect -682 367 -666 401
rect -632 367 -616 401
rect -682 351 -616 367
rect -564 401 -498 417
rect -564 367 -548 401
rect -514 367 -498 401
rect -564 351 -498 367
rect -446 401 -380 417
rect -446 367 -430 401
rect -396 367 -380 401
rect -446 351 -380 367
rect -328 401 -262 417
rect -328 367 -312 401
rect -278 367 -262 401
rect -328 351 -262 367
rect -210 401 -144 417
rect -210 367 -194 401
rect -160 367 -144 401
rect -210 351 -144 367
rect -92 401 -26 417
rect -92 367 -76 401
rect -42 367 -26 401
rect -92 351 -26 367
rect 26 401 92 417
rect 26 367 42 401
rect 76 367 92 401
rect 26 351 92 367
rect 144 401 210 417
rect 144 367 160 401
rect 194 367 210 401
rect 144 351 210 367
rect 262 401 328 417
rect 262 367 278 401
rect 312 367 328 401
rect 262 351 328 367
rect 380 401 446 417
rect 380 367 396 401
rect 430 367 446 401
rect 380 351 446 367
rect 498 401 564 417
rect 498 367 514 401
rect 548 367 564 401
rect 498 351 564 367
rect 616 401 682 417
rect 616 367 632 401
rect 666 367 682 401
rect 616 351 682 367
rect -679 329 -619 351
rect -561 329 -501 351
rect -443 329 -383 351
rect -325 329 -265 351
rect -207 329 -147 351
rect -89 329 -29 351
rect 29 329 89 351
rect 147 329 207 351
rect 265 329 325 351
rect 383 329 443 351
rect 501 329 561 351
rect 619 329 679 351
rect -679 -417 -619 -391
rect -561 -417 -501 -391
rect -443 -417 -383 -391
rect -325 -417 -265 -391
rect -207 -417 -147 -391
rect -89 -417 -29 -391
rect 29 -417 89 -391
rect 147 -417 207 -391
rect 265 -417 325 -391
rect 383 -417 443 -391
rect 501 -417 561 -391
rect 619 -417 679 -391
<< polycont >>
rect -666 367 -632 401
rect -548 367 -514 401
rect -430 367 -396 401
rect -312 367 -278 401
rect -194 367 -160 401
rect -76 367 -42 401
rect 42 367 76 401
rect 160 367 194 401
rect 278 367 312 401
rect 396 367 430 401
rect 514 367 548 401
rect 632 367 666 401
<< locali >>
rect -839 469 -743 503
rect 743 469 839 503
rect -839 407 -805 469
rect 805 407 839 469
rect -682 367 -666 401
rect -632 367 -616 401
rect -564 367 -548 401
rect -514 367 -498 401
rect -446 367 -430 401
rect -396 367 -380 401
rect -328 367 -312 401
rect -278 367 -262 401
rect -210 367 -194 401
rect -160 367 -144 401
rect -92 367 -76 401
rect -42 367 -26 401
rect 26 367 42 401
rect 76 367 92 401
rect 144 367 160 401
rect 194 367 210 401
rect 262 367 278 401
rect 312 367 328 401
rect 380 367 396 401
rect 430 367 446 401
rect 498 367 514 401
rect 548 367 564 401
rect 616 367 632 401
rect 666 367 682 401
rect -725 317 -691 333
rect -725 -395 -691 -379
rect -607 317 -573 333
rect -607 -395 -573 -379
rect -489 317 -455 333
rect -489 -395 -455 -379
rect -371 317 -337 333
rect -371 -395 -337 -379
rect -253 317 -219 333
rect -253 -395 -219 -379
rect -135 317 -101 333
rect -135 -395 -101 -379
rect -17 317 17 333
rect -17 -395 17 -379
rect 101 317 135 333
rect 101 -395 135 -379
rect 219 317 253 333
rect 219 -395 253 -379
rect 337 317 371 333
rect 337 -395 371 -379
rect 455 317 489 333
rect 455 -395 489 -379
rect 573 317 607 333
rect 573 -395 607 -379
rect 691 317 725 333
rect 691 -395 725 -379
rect -839 -469 -805 -407
rect 805 -469 839 -407
rect -839 -503 -743 -469
rect 743 -503 839 -469
<< viali >>
rect -666 367 -632 401
rect -548 367 -514 401
rect -430 367 -396 401
rect -312 367 -278 401
rect -194 367 -160 401
rect -76 367 -42 401
rect 42 367 76 401
rect 160 367 194 401
rect 278 367 312 401
rect 396 367 430 401
rect 514 367 548 401
rect 632 367 666 401
rect -725 -379 -691 317
rect -607 -379 -573 317
rect -489 -379 -455 317
rect -371 -379 -337 317
rect -253 -379 -219 317
rect -135 -379 -101 317
rect -17 -379 17 317
rect 101 -379 135 317
rect 219 -379 253 317
rect 337 -379 371 317
rect 455 -379 489 317
rect 573 -379 607 317
rect 691 -379 725 317
<< metal1 >>
rect -678 401 -620 407
rect -678 367 -666 401
rect -632 367 -620 401
rect -678 361 -620 367
rect -560 401 -502 407
rect -560 367 -548 401
rect -514 367 -502 401
rect -560 361 -502 367
rect -442 401 -384 407
rect -442 367 -430 401
rect -396 367 -384 401
rect -442 361 -384 367
rect -324 401 -266 407
rect -324 367 -312 401
rect -278 367 -266 401
rect -324 361 -266 367
rect -206 401 -148 407
rect -206 367 -194 401
rect -160 367 -148 401
rect -206 361 -148 367
rect -88 401 -30 407
rect -88 367 -76 401
rect -42 367 -30 401
rect -88 361 -30 367
rect 30 401 88 407
rect 30 367 42 401
rect 76 367 88 401
rect 30 361 88 367
rect 148 401 206 407
rect 148 367 160 401
rect 194 367 206 401
rect 148 361 206 367
rect 266 401 324 407
rect 266 367 278 401
rect 312 367 324 401
rect 266 361 324 367
rect 384 401 442 407
rect 384 367 396 401
rect 430 367 442 401
rect 384 361 442 367
rect 502 401 560 407
rect 502 367 514 401
rect 548 367 560 401
rect 502 361 560 367
rect 620 401 678 407
rect 620 367 632 401
rect 666 367 678 401
rect 620 361 678 367
rect -731 317 -685 329
rect -731 -379 -725 317
rect -691 -379 -685 317
rect -731 -391 -685 -379
rect -613 317 -567 329
rect -613 -379 -607 317
rect -573 -379 -567 317
rect -613 -391 -567 -379
rect -495 317 -449 329
rect -495 -379 -489 317
rect -455 -379 -449 317
rect -495 -391 -449 -379
rect -377 317 -331 329
rect -377 -379 -371 317
rect -337 -379 -331 317
rect -377 -391 -331 -379
rect -259 317 -213 329
rect -259 -379 -253 317
rect -219 -379 -213 317
rect -259 -391 -213 -379
rect -141 317 -95 329
rect -141 -379 -135 317
rect -101 -379 -95 317
rect -141 -391 -95 -379
rect -23 317 23 329
rect -23 -379 -17 317
rect 17 -379 23 317
rect -23 -391 23 -379
rect 95 317 141 329
rect 95 -379 101 317
rect 135 -379 141 317
rect 95 -391 141 -379
rect 213 317 259 329
rect 213 -379 219 317
rect 253 -379 259 317
rect 213 -391 259 -379
rect 331 317 377 329
rect 331 -379 337 317
rect 371 -379 377 317
rect 331 -391 377 -379
rect 449 317 495 329
rect 449 -379 455 317
rect 489 -379 495 317
rect 449 -391 495 -379
rect 567 317 613 329
rect 567 -379 573 317
rect 607 -379 613 317
rect 567 -391 613 -379
rect 685 317 731 329
rect 685 -379 691 317
rect 725 -379 731 317
rect 685 -391 731 -379
<< labels >>
flabel metal1 -649 384 -649 384 0 FreeSans 240 0 0 0 G
flabel metal1 -531 384 -531 384 0 FreeSans 240 0 0 0 G
flabel metal1 -413 384 -413 384 0 FreeSans 240 0 0 0 G
flabel metal1 -295 384 -295 384 0 FreeSans 240 0 0 0 G
flabel metal1 -177 384 -177 384 0 FreeSans 240 0 0 0 G
flabel metal1 -59 384 -59 384 0 FreeSans 240 0 0 0 G
flabel metal1 59 384 59 384 0 FreeSans 240 0 0 0 G
flabel metal1 177 384 177 384 0 FreeSans 240 0 0 0 G
flabel metal1 295 384 295 384 0 FreeSans 240 0 0 0 G
flabel metal1 413 384 413 384 0 FreeSans 240 0 0 0 G
flabel metal1 531 384 531 384 0 FreeSans 240 0 0 0 G
flabel metal1 649 384 649 384 0 FreeSans 240 0 0 0 G
flabel metal1 -708 -31 -708 -31 0 FreeSans 240 0 0 0 D
flabel metal1 -590 -31 -590 -31 0 FreeSans 240 0 0 0 S
flabel metal1 -472 -31 -472 -31 0 FreeSans 240 0 0 0 D
flabel metal1 -354 -31 -354 -31 0 FreeSans 240 0 0 0 S
flabel metal1 -236 -31 -236 -31 0 FreeSans 240 0 0 0 D
flabel metal1 -118 -31 -118 -31 0 FreeSans 240 0 0 0 S
flabel metal1 0 -31 0 -31 0 FreeSans 240 0 0 0 D
flabel metal1 118 -31 118 -31 0 FreeSans 240 0 0 0 S
flabel metal1 236 -31 236 -31 0 FreeSans 240 0 0 0 D
flabel metal1 354 -31 354 -31 0 FreeSans 240 0 0 0 S
flabel metal1 472 -31 472 -31 0 FreeSans 240 0 0 0 D
flabel metal1 590 -31 590 -31 0 FreeSans 240 0 0 0 S
flabel metal1 708 -31 708 -31 0 FreeSans 240 0 0 0 D
<< properties >>
string FIXED_BBOX -822 -486 822 486
<< end >>

