magic
tech sky130A
magscale 1 2
timestamp 1679988684
<< checkpaint >>
rect -1210 4810 11410 4860
rect -1260 -1210 11460 4810
rect -1260 -1260 11410 -1210
<< viali >>
rect 1144 3078 1178 3112
rect 3420 3078 3454 3112
rect 3944 3078 3978 3112
rect 6220 3078 6254 3112
rect 6744 3078 6778 3112
rect 9020 3078 9054 3112
rect 1144 3006 1178 3040
rect 3420 3006 3454 3040
rect 3944 3006 3978 3040
rect 6220 3006 6254 3040
rect 6744 3006 6778 3040
rect 9020 3006 9054 3040
rect 1144 2934 1178 2968
rect 3420 2934 3454 2968
rect 3944 2934 3978 2968
rect 6220 2934 6254 2968
rect 6744 2934 6778 2968
rect 9020 2934 9054 2968
rect 1144 2862 1178 2896
rect 3420 2862 3454 2896
rect 3944 2862 3978 2896
rect 6220 2862 6254 2896
rect 6744 2862 6778 2896
rect 9020 2862 9054 2896
rect 1144 2790 1178 2824
rect 3420 2790 3454 2824
rect 3944 2790 3978 2824
rect 6220 2790 6254 2824
rect 6744 2790 6778 2824
rect 9020 2790 9054 2824
rect 1144 2718 1178 2752
rect 3420 2718 3454 2752
rect 3944 2718 3978 2752
rect 6220 2718 6254 2752
rect 6744 2718 6778 2752
rect 9020 2718 9054 2752
rect 278 2618 312 2652
rect 688 2618 722 2652
rect 1144 2646 1178 2680
rect 3420 2646 3454 2680
rect 3944 2646 3978 2680
rect 6220 2646 6254 2680
rect 6744 2646 6778 2680
rect 9020 2646 9054 2680
rect 9478 2618 9512 2652
rect 9888 2618 9922 2652
rect 278 2546 312 2580
rect 688 2546 722 2580
rect 1144 2574 1178 2608
rect 3420 2574 3454 2608
rect 3944 2574 3978 2608
rect 6220 2574 6254 2608
rect 6744 2574 6778 2608
rect 9020 2574 9054 2608
rect 9478 2546 9512 2580
rect 9888 2546 9922 2580
rect 278 2474 312 2508
rect 688 2474 722 2508
rect 1144 2502 1178 2536
rect 3420 2502 3454 2536
rect 3944 2502 3978 2536
rect 6220 2502 6254 2536
rect 6744 2502 6778 2536
rect 9020 2502 9054 2536
rect 9478 2474 9512 2508
rect 9888 2474 9922 2508
rect 278 2402 312 2436
rect 688 2402 722 2436
rect 1144 2430 1178 2464
rect 3420 2430 3454 2464
rect 3944 2430 3978 2464
rect 6220 2430 6254 2464
rect 6744 2430 6778 2464
rect 9020 2430 9054 2464
rect 9478 2402 9512 2436
rect 9888 2402 9922 2436
rect 278 2330 312 2364
rect 688 2330 722 2364
rect 1144 2358 1178 2392
rect 3420 2358 3454 2392
rect 3944 2358 3978 2392
rect 6220 2358 6254 2392
rect 6744 2358 6778 2392
rect 9020 2358 9054 2392
rect 9478 2330 9512 2364
rect 9888 2330 9922 2364
rect 278 2258 312 2292
rect 688 2258 722 2292
rect 1144 2286 1178 2320
rect 3420 2286 3454 2320
rect 3944 2286 3978 2320
rect 6220 2286 6254 2320
rect 6744 2286 6778 2320
rect 9020 2286 9054 2320
rect 9478 2258 9512 2292
rect 9888 2258 9922 2292
rect 278 2186 312 2220
rect 688 2186 722 2220
rect 9478 2186 9512 2220
rect 9888 2186 9922 2220
rect 278 2114 312 2148
rect 688 2114 722 2148
rect 9478 2114 9512 2148
rect 9888 2114 9922 2148
rect 278 2042 312 2076
rect 688 2042 722 2076
rect 9478 2042 9512 2076
rect 9888 2042 9922 2076
rect 278 1970 312 2004
rect 688 1970 722 2004
rect 9478 1970 9512 2004
rect 9888 1970 9922 2004
rect 278 1898 312 1932
rect 688 1898 722 1932
rect 9478 1898 9512 1932
rect 9888 1898 9922 1932
rect 278 1826 312 1860
rect 688 1826 722 1860
rect 9478 1826 9512 1860
rect 9888 1826 9922 1860
rect 278 1754 312 1788
rect 688 1754 722 1788
rect 9478 1754 9512 1788
rect 9888 1754 9922 1788
rect 278 1682 312 1716
rect 688 1682 722 1716
rect 9478 1682 9512 1716
rect 9888 1682 9922 1716
rect 278 1610 312 1644
rect 688 1610 722 1644
rect 9478 1610 9512 1644
rect 9888 1610 9922 1644
rect 278 1538 312 1572
rect 688 1538 722 1572
rect 9478 1538 9512 1572
rect 9888 1538 9922 1572
rect 278 1466 312 1500
rect 688 1466 722 1500
rect 9478 1466 9512 1500
rect 9888 1466 9922 1500
rect 278 1394 312 1428
rect 688 1394 722 1428
rect 9478 1394 9512 1428
rect 9888 1394 9922 1428
rect 278 1322 312 1356
rect 688 1322 722 1356
rect 9478 1322 9512 1356
rect 9888 1322 9922 1356
rect 278 1250 312 1284
rect 688 1250 722 1284
rect 1144 1278 1178 1312
rect 3420 1278 3454 1312
rect 3944 1278 3978 1312
rect 6220 1278 6254 1312
rect 6744 1278 6778 1312
rect 9020 1278 9054 1312
rect 9478 1250 9512 1284
rect 9888 1250 9922 1284
rect 278 1178 312 1212
rect 688 1178 722 1212
rect 1144 1206 1178 1240
rect 3420 1206 3454 1240
rect 3944 1206 3978 1240
rect 6220 1206 6254 1240
rect 6744 1206 6778 1240
rect 9020 1206 9054 1240
rect 9478 1178 9512 1212
rect 9888 1178 9922 1212
rect 278 1106 312 1140
rect 688 1106 722 1140
rect 1144 1134 1178 1168
rect 3420 1134 3454 1168
rect 3944 1134 3978 1168
rect 6220 1134 6254 1168
rect 6744 1134 6778 1168
rect 9020 1134 9054 1168
rect 9478 1106 9512 1140
rect 9888 1106 9922 1140
rect 278 1034 312 1068
rect 688 1034 722 1068
rect 1144 1062 1178 1096
rect 3420 1062 3454 1096
rect 3944 1062 3978 1096
rect 6220 1062 6254 1096
rect 6744 1062 6778 1096
rect 9020 1062 9054 1096
rect 9478 1034 9512 1068
rect 9888 1034 9922 1068
rect 278 962 312 996
rect 688 962 722 996
rect 1144 990 1178 1024
rect 3420 990 3454 1024
rect 3944 990 3978 1024
rect 6220 990 6254 1024
rect 6744 990 6778 1024
rect 9020 990 9054 1024
rect 9478 962 9512 996
rect 9888 962 9922 996
rect 278 890 312 924
rect 688 890 722 924
rect 1144 918 1178 952
rect 3420 918 3454 952
rect 3944 918 3978 952
rect 6220 918 6254 952
rect 6744 918 6778 952
rect 9020 918 9054 952
rect 9478 890 9512 924
rect 9888 890 9922 924
rect 278 818 312 852
rect 688 818 722 852
rect 1144 846 1178 880
rect 3420 846 3454 880
rect 3944 846 3978 880
rect 6220 846 6254 880
rect 6744 846 6778 880
rect 9020 846 9054 880
rect 9478 818 9512 852
rect 9888 818 9922 852
rect 278 746 312 780
rect 688 746 722 780
rect 1144 774 1178 808
rect 3420 774 3454 808
rect 3944 774 3978 808
rect 6220 774 6254 808
rect 6744 774 6778 808
rect 9020 774 9054 808
rect 9478 746 9512 780
rect 9888 746 9922 780
rect 1144 702 1178 736
rect 3420 702 3454 736
rect 3944 702 3978 736
rect 6220 702 6254 736
rect 6744 702 6778 736
rect 9020 702 9054 736
rect 1144 630 1178 664
rect 3420 630 3454 664
rect 3944 630 3978 664
rect 6220 630 6254 664
rect 6744 630 6778 664
rect 9020 630 9054 664
rect 1144 558 1178 592
rect 3420 558 3454 592
rect 3944 558 3978 592
rect 6220 558 6254 592
rect 6744 558 6778 592
rect 9020 558 9054 592
rect 1144 486 1178 520
rect 3420 486 3454 520
rect 3944 486 3978 520
rect 6220 486 6254 520
rect 6744 486 6778 520
rect 9020 486 9054 520
<< metal1 >>
rect 50 3550 150 3600
rect 250 3550 350 3600
rect 450 3550 550 3600
rect 650 3550 750 3600
rect 850 3550 950 3600
rect 1050 3550 1150 3600
rect 1250 3550 1350 3600
rect 1450 3550 1550 3600
rect 1650 3550 1750 3600
rect 1850 3550 1950 3600
rect 2050 3550 2150 3600
rect 2250 3550 2350 3600
rect 2450 3550 2550 3600
rect 2650 3550 2750 3600
rect 2850 3550 2950 3600
rect 3050 3550 3150 3600
rect 3250 3550 3350 3600
rect 3450 3550 3550 3600
rect 3650 3550 3750 3600
rect 3850 3550 3950 3600
rect 4050 3550 4150 3600
rect 4250 3550 4350 3600
rect 4450 3550 4550 3600
rect 4650 3550 4750 3600
rect 4850 3550 4950 3600
rect 5050 3550 5150 3600
rect 5250 3550 5350 3600
rect 5450 3550 5550 3600
rect 5650 3550 5750 3600
rect 5850 3550 5950 3600
rect 6050 3550 6150 3600
rect 6250 3550 6350 3600
rect 6450 3550 6550 3600
rect 6650 3550 6750 3600
rect 6850 3550 6950 3600
rect 7050 3550 7150 3600
rect 7250 3550 7350 3600
rect 7450 3550 7550 3600
rect 7650 3550 7750 3600
rect 7850 3550 7950 3600
rect 8050 3550 8150 3600
rect 8250 3550 8350 3600
rect 8450 3550 8550 3600
rect 8650 3550 8750 3600
rect 8850 3550 8950 3600
rect 9050 3550 9150 3600
rect 9250 3550 9350 3600
rect 9450 3550 9550 3600
rect 9650 3550 9750 3600
rect 9850 3550 9950 3600
rect 10050 3550 10150 3600
rect 0 3450 10200 3550
rect 50 3350 150 3450
rect 250 3350 350 3450
rect 450 3350 550 3450
rect 650 3350 750 3450
rect 850 3350 950 3450
rect 1050 3400 1150 3450
rect 1250 3400 1350 3450
rect 1450 3400 1550 3450
rect 1650 3400 1750 3450
rect 1850 3400 1950 3450
rect 2050 3400 2150 3450
rect 2250 3400 2350 3450
rect 2450 3400 2550 3450
rect 2650 3400 2750 3450
rect 2850 3400 2950 3450
rect 3050 3400 3150 3450
rect 3250 3400 3350 3450
rect 3450 3400 3550 3450
rect 3650 3350 3750 3450
rect 3850 3400 3950 3450
rect 4050 3400 4150 3450
rect 4250 3400 4350 3450
rect 4450 3400 4550 3450
rect 4650 3400 4750 3450
rect 4850 3400 4950 3450
rect 5050 3400 5150 3450
rect 5250 3400 5350 3450
rect 5450 3400 5550 3450
rect 5650 3400 5750 3450
rect 5850 3400 5950 3450
rect 6050 3400 6150 3450
rect 6250 3400 6350 3450
rect 6450 3350 6550 3450
rect 6650 3400 6750 3450
rect 6850 3400 6950 3450
rect 7050 3400 7150 3450
rect 7250 3400 7350 3450
rect 7450 3400 7550 3450
rect 7650 3400 7750 3450
rect 7850 3400 7950 3450
rect 8050 3400 8150 3450
rect 8250 3400 8350 3450
rect 8450 3400 8550 3450
rect 8650 3400 8750 3450
rect 8850 3400 8950 3450
rect 9050 3400 9150 3450
rect 9250 3350 9350 3450
rect 9450 3350 9550 3450
rect 9650 3350 9750 3450
rect 9850 3350 9950 3450
rect 10050 3350 10150 3450
rect 0 3250 1000 3350
rect 3600 3250 3800 3350
rect 6400 3250 6600 3350
rect 9200 3250 10200 3350
rect 50 3150 150 3250
rect 250 3150 350 3250
rect 450 3150 550 3250
rect 650 3150 750 3250
rect 850 3150 950 3250
rect 0 3050 1000 3150
rect 1122 3112 1202 3158
rect 1122 3078 1144 3112
rect 1178 3078 1202 3112
rect 50 2950 150 3050
rect 250 3000 350 3050
rect 0 2850 200 2950
rect 50 2750 150 2850
rect 0 2650 200 2750
rect 254 2652 334 2690
rect 50 2550 150 2650
rect 254 2618 278 2652
rect 312 2618 334 2652
rect 450 2650 550 3050
rect 650 3000 750 3050
rect 850 2950 950 3050
rect 1122 3040 1202 3078
rect 1122 3006 1144 3040
rect 1178 3006 1202 3040
rect 1122 2968 1202 3006
rect 800 2850 1000 2950
rect 1122 2934 1144 2968
rect 1178 2934 1202 2968
rect 1122 2896 1202 2934
rect 1122 2862 1144 2896
rect 1178 2862 1202 2896
rect 850 2750 950 2850
rect 1122 2824 1202 2862
rect 1122 2790 1144 2824
rect 1178 2790 1202 2824
rect 1122 2752 1202 2790
rect 664 2652 744 2690
rect 254 2580 334 2618
rect 254 2550 278 2580
rect 0 2546 278 2550
rect 312 2546 334 2580
rect 0 2508 334 2546
rect 0 2474 278 2508
rect 312 2474 334 2508
rect 0 2450 334 2474
rect 50 2350 150 2450
rect 254 2436 334 2450
rect 254 2402 278 2436
rect 312 2402 334 2436
rect 254 2364 334 2402
rect 254 2350 278 2364
rect 0 2330 278 2350
rect 312 2330 334 2364
rect 0 2292 334 2330
rect 0 2258 278 2292
rect 312 2258 334 2292
rect 0 2250 334 2258
rect 50 2150 150 2250
rect 254 2220 334 2250
rect 254 2186 278 2220
rect 312 2186 334 2220
rect 254 2150 334 2186
rect 0 2148 334 2150
rect 0 2114 278 2148
rect 312 2114 334 2148
rect 0 2076 334 2114
rect 0 2050 278 2076
rect 50 1950 150 2050
rect 254 2042 278 2050
rect 312 2042 334 2076
rect 254 2004 334 2042
rect 254 1970 278 2004
rect 312 1970 334 2004
rect 254 1950 334 1970
rect 0 1932 334 1950
rect 0 1898 278 1932
rect 312 1898 334 1932
rect 0 1860 334 1898
rect 0 1850 278 1860
rect 50 1750 150 1850
rect 254 1826 278 1850
rect 312 1826 334 1860
rect 254 1788 334 1826
rect 254 1754 278 1788
rect 312 1754 334 1788
rect 254 1750 334 1754
rect 0 1716 334 1750
rect 0 1682 278 1716
rect 312 1682 334 1716
rect 0 1650 334 1682
rect 50 1550 150 1650
rect 254 1644 334 1650
rect 254 1610 278 1644
rect 312 1610 334 1644
rect 254 1572 334 1610
rect 254 1550 278 1572
rect 0 1538 278 1550
rect 312 1538 334 1572
rect 0 1500 334 1538
rect 0 1466 278 1500
rect 312 1466 334 1500
rect 0 1450 334 1466
rect 50 1350 150 1450
rect 254 1428 334 1450
rect 254 1394 278 1428
rect 312 1394 334 1428
rect 254 1356 334 1394
rect 254 1350 278 1356
rect 0 1322 278 1350
rect 312 1322 334 1356
rect 0 1284 334 1322
rect 0 1250 278 1284
rect 312 1250 334 1284
rect 50 1150 150 1250
rect 254 1212 334 1250
rect 254 1178 278 1212
rect 312 1178 334 1212
rect 254 1150 334 1178
rect 0 1140 334 1150
rect 0 1106 278 1140
rect 312 1106 334 1140
rect 0 1068 334 1106
rect 0 1050 278 1068
rect 50 950 150 1050
rect 254 1034 278 1050
rect 312 1034 334 1068
rect 254 996 334 1034
rect 254 962 278 996
rect 312 962 334 996
rect 254 950 334 962
rect 0 924 334 950
rect 0 890 278 924
rect 312 890 334 924
rect 0 852 334 890
rect 0 850 278 852
rect 50 750 150 850
rect 254 818 278 850
rect 312 818 334 852
rect 254 780 334 818
rect 0 650 200 750
rect 254 746 278 780
rect 312 746 334 780
rect 254 708 334 746
rect 664 2618 688 2652
rect 722 2618 744 2652
rect 800 2650 1000 2750
rect 1122 2718 1144 2752
rect 1178 2718 1202 2752
rect 1122 2680 1202 2718
rect 664 2580 744 2618
rect 664 2546 688 2580
rect 722 2550 744 2580
rect 850 2550 950 2650
rect 1122 2646 1144 2680
rect 1178 2646 1202 2680
rect 1122 2608 1202 2646
rect 1122 2574 1144 2608
rect 1178 2574 1202 2608
rect 722 2546 1000 2550
rect 664 2508 1000 2546
rect 664 2474 688 2508
rect 722 2474 1000 2508
rect 664 2450 1000 2474
rect 1122 2536 1202 2574
rect 1122 2502 1144 2536
rect 1178 2502 1202 2536
rect 1122 2464 1202 2502
rect 664 2436 744 2450
rect 664 2402 688 2436
rect 722 2402 744 2436
rect 664 2364 744 2402
rect 664 2330 688 2364
rect 722 2350 744 2364
rect 850 2350 950 2450
rect 1122 2430 1144 2464
rect 1178 2430 1202 2464
rect 1122 2392 1202 2430
rect 1122 2358 1144 2392
rect 1178 2358 1202 2392
rect 722 2330 1000 2350
rect 664 2292 1000 2330
rect 664 2258 688 2292
rect 722 2258 1000 2292
rect 664 2250 1000 2258
rect 1122 2320 1202 2358
rect 1122 2286 1144 2320
rect 1178 2286 1202 2320
rect 664 2220 744 2250
rect 664 2186 688 2220
rect 722 2186 744 2220
rect 664 2150 744 2186
rect 850 2150 950 2250
rect 1122 2240 1202 2286
rect 3398 3112 3478 3158
rect 3650 3150 3750 3250
rect 3398 3078 3420 3112
rect 3454 3078 3478 3112
rect 3398 3040 3478 3078
rect 3600 3050 3800 3150
rect 3922 3112 4000 3158
rect 3922 3078 3944 3112
rect 3978 3078 4000 3112
rect 3398 3006 3420 3040
rect 3454 3006 3478 3040
rect 3398 2968 3478 3006
rect 3398 2934 3420 2968
rect 3454 2934 3478 2968
rect 3650 2950 3750 3050
rect 3922 3040 4000 3078
rect 3922 3006 3944 3040
rect 3978 3006 4000 3040
rect 3922 2968 4000 3006
rect 3398 2896 3478 2934
rect 3398 2862 3420 2896
rect 3454 2862 3478 2896
rect 3398 2824 3478 2862
rect 3600 2850 3800 2950
rect 3922 2934 3944 2968
rect 3978 2934 4000 2968
rect 3922 2896 4000 2934
rect 3922 2862 3944 2896
rect 3978 2862 4000 2896
rect 3398 2790 3420 2824
rect 3454 2790 3478 2824
rect 3398 2752 3478 2790
rect 3398 2718 3420 2752
rect 3454 2718 3478 2752
rect 3650 2750 3750 2850
rect 3922 2824 4000 2862
rect 3922 2790 3944 2824
rect 3978 2790 4000 2824
rect 3922 2752 4000 2790
rect 3398 2680 3478 2718
rect 3398 2646 3420 2680
rect 3454 2646 3478 2680
rect 3600 2650 3800 2750
rect 3922 2718 3944 2752
rect 3978 2718 4000 2752
rect 3922 2680 4000 2718
rect 3398 2608 3478 2646
rect 3398 2574 3420 2608
rect 3454 2574 3478 2608
rect 3398 2536 3478 2574
rect 3650 2550 3750 2650
rect 3922 2646 3944 2680
rect 3978 2646 4000 2680
rect 3922 2608 4000 2646
rect 3922 2574 3944 2608
rect 3978 2574 4000 2608
rect 3398 2502 3420 2536
rect 3454 2502 3478 2536
rect 3398 2464 3478 2502
rect 3398 2430 3420 2464
rect 3454 2430 3478 2464
rect 3600 2450 3800 2550
rect 3922 2536 4000 2574
rect 3922 2502 3944 2536
rect 3978 2502 4000 2536
rect 3922 2464 4000 2502
rect 3398 2392 3478 2430
rect 3398 2358 3420 2392
rect 3454 2358 3478 2392
rect 3398 2320 3478 2358
rect 3650 2350 3750 2450
rect 3922 2430 3944 2464
rect 3978 2430 4000 2464
rect 3922 2392 4000 2430
rect 3922 2358 3944 2392
rect 3978 2358 4000 2392
rect 3398 2286 3420 2320
rect 3454 2286 3478 2320
rect 3398 2240 3478 2286
rect 3600 2250 3800 2350
rect 3922 2320 4000 2358
rect 3922 2286 3944 2320
rect 3978 2286 4000 2320
rect 3650 2150 3750 2250
rect 3922 2240 4000 2286
rect 6198 3112 6278 3158
rect 6450 3150 6550 3250
rect 6198 3078 6220 3112
rect 6254 3078 6278 3112
rect 6198 3040 6278 3078
rect 6400 3050 6600 3150
rect 6722 3112 6802 3158
rect 6722 3078 6744 3112
rect 6778 3078 6802 3112
rect 6198 3006 6220 3040
rect 6254 3006 6278 3040
rect 6198 2968 6278 3006
rect 6198 2934 6220 2968
rect 6254 2934 6278 2968
rect 6450 2950 6550 3050
rect 6722 3040 6802 3078
rect 6722 3006 6744 3040
rect 6778 3006 6802 3040
rect 6722 2968 6802 3006
rect 6198 2896 6278 2934
rect 6198 2862 6220 2896
rect 6254 2862 6278 2896
rect 6198 2824 6278 2862
rect 6400 2850 6600 2950
rect 6722 2934 6744 2968
rect 6778 2934 6802 2968
rect 6722 2896 6802 2934
rect 6722 2862 6744 2896
rect 6778 2862 6802 2896
rect 6198 2790 6220 2824
rect 6254 2790 6278 2824
rect 6198 2752 6278 2790
rect 6198 2718 6220 2752
rect 6254 2718 6278 2752
rect 6450 2750 6550 2850
rect 6722 2824 6802 2862
rect 6722 2790 6744 2824
rect 6778 2790 6802 2824
rect 6722 2752 6802 2790
rect 6198 2680 6278 2718
rect 6198 2646 6220 2680
rect 6254 2646 6278 2680
rect 6400 2650 6600 2750
rect 6722 2718 6744 2752
rect 6778 2718 6802 2752
rect 6722 2680 6802 2718
rect 6198 2608 6278 2646
rect 6198 2574 6220 2608
rect 6254 2574 6278 2608
rect 6198 2536 6278 2574
rect 6450 2550 6550 2650
rect 6722 2646 6744 2680
rect 6778 2646 6802 2680
rect 6722 2608 6802 2646
rect 6722 2574 6744 2608
rect 6778 2574 6802 2608
rect 6198 2502 6220 2536
rect 6254 2502 6278 2536
rect 6198 2464 6278 2502
rect 6198 2430 6220 2464
rect 6254 2430 6278 2464
rect 6400 2450 6600 2550
rect 6722 2536 6802 2574
rect 6722 2502 6744 2536
rect 6778 2502 6802 2536
rect 6722 2464 6802 2502
rect 6198 2392 6278 2430
rect 6198 2358 6220 2392
rect 6254 2358 6278 2392
rect 6198 2320 6278 2358
rect 6450 2350 6550 2450
rect 6722 2430 6744 2464
rect 6778 2430 6802 2464
rect 6722 2392 6802 2430
rect 6722 2358 6744 2392
rect 6778 2358 6802 2392
rect 6198 2286 6220 2320
rect 6254 2286 6278 2320
rect 6198 2240 6278 2286
rect 6400 2250 6600 2350
rect 6722 2320 6802 2358
rect 6722 2286 6744 2320
rect 6778 2286 6802 2320
rect 6450 2150 6550 2250
rect 6722 2240 6802 2286
rect 8996 3112 9078 3158
rect 9250 3150 9350 3250
rect 9450 3150 9550 3250
rect 9650 3150 9750 3250
rect 9850 3150 9950 3250
rect 10050 3150 10150 3250
rect 8996 3078 9020 3112
rect 9054 3078 9078 3112
rect 8996 3040 9078 3078
rect 9200 3050 10200 3150
rect 8996 3006 9020 3040
rect 9054 3006 9078 3040
rect 8996 2968 9078 3006
rect 8996 2934 9020 2968
rect 9054 2934 9078 2968
rect 9250 2950 9350 3050
rect 9450 3000 9550 3050
rect 8996 2896 9078 2934
rect 8996 2862 9020 2896
rect 9054 2862 9078 2896
rect 8996 2824 9078 2862
rect 9200 2850 9400 2950
rect 8996 2790 9020 2824
rect 9054 2790 9078 2824
rect 8996 2752 9078 2790
rect 8996 2718 9020 2752
rect 9054 2718 9078 2752
rect 9250 2750 9350 2850
rect 8996 2680 9078 2718
rect 8996 2646 9020 2680
rect 9054 2646 9078 2680
rect 9200 2650 9400 2750
rect 9454 2652 9534 2690
rect 8996 2608 9078 2646
rect 8996 2574 9020 2608
rect 9054 2574 9078 2608
rect 8996 2536 9078 2574
rect 9250 2550 9350 2650
rect 9454 2618 9478 2652
rect 9512 2618 9534 2652
rect 9650 2650 9750 3050
rect 9850 3000 9950 3050
rect 10050 2950 10150 3050
rect 10000 2850 10200 2950
rect 10050 2750 10150 2850
rect 9864 2652 9944 2690
rect 9454 2580 9534 2618
rect 9454 2550 9478 2580
rect 8996 2502 9020 2536
rect 9054 2502 9078 2536
rect 8996 2464 9078 2502
rect 8996 2430 9020 2464
rect 9054 2430 9078 2464
rect 9200 2546 9478 2550
rect 9512 2546 9534 2580
rect 9200 2508 9534 2546
rect 9200 2474 9478 2508
rect 9512 2474 9534 2508
rect 9200 2450 9534 2474
rect 8996 2392 9078 2430
rect 8996 2358 9020 2392
rect 9054 2358 9078 2392
rect 8996 2320 9078 2358
rect 9250 2350 9350 2450
rect 9454 2436 9534 2450
rect 9454 2402 9478 2436
rect 9512 2402 9534 2436
rect 9454 2364 9534 2402
rect 9454 2350 9478 2364
rect 8996 2286 9020 2320
rect 9054 2286 9078 2320
rect 8996 2240 9078 2286
rect 9200 2330 9478 2350
rect 9512 2330 9534 2364
rect 9200 2292 9534 2330
rect 9200 2258 9478 2292
rect 9512 2258 9534 2292
rect 9200 2250 9534 2258
rect 9250 2150 9350 2250
rect 9454 2220 9534 2250
rect 9454 2186 9478 2220
rect 9512 2186 9534 2220
rect 9454 2150 9534 2186
rect 664 2148 1000 2150
rect 664 2114 688 2148
rect 722 2114 1000 2148
rect 664 2076 1000 2114
rect 664 2042 688 2076
rect 722 2050 1000 2076
rect 3600 2050 3800 2150
rect 6400 2050 6600 2150
rect 9200 2148 9534 2150
rect 9200 2114 9478 2148
rect 9512 2114 9534 2148
rect 9200 2076 9534 2114
rect 9200 2050 9478 2076
rect 722 2042 744 2050
rect 664 2004 744 2042
rect 664 1970 688 2004
rect 722 1970 744 2004
rect 664 1950 744 1970
rect 850 1950 950 2050
rect 1050 1950 1150 2000
rect 1250 1950 1350 2000
rect 1450 1950 1550 2000
rect 1650 1950 1750 2000
rect 1850 1950 1950 2000
rect 2050 1950 2150 2000
rect 2250 1950 2350 2000
rect 2450 1950 2550 2000
rect 2650 1950 2750 2000
rect 2850 1950 2950 2000
rect 3050 1950 3150 2000
rect 3250 1950 3350 2000
rect 3450 1950 3550 2000
rect 3650 1950 3750 2050
rect 3850 1950 3950 2000
rect 4050 1950 4150 2000
rect 4250 1950 4350 2000
rect 4450 1950 4550 2000
rect 4650 1950 4750 2000
rect 4850 1950 4950 2000
rect 5050 1950 5150 2000
rect 5250 1950 5350 2000
rect 5450 1950 5550 2000
rect 5650 1950 5750 2000
rect 5850 1950 5950 2000
rect 6050 1950 6150 2000
rect 6250 1950 6350 2000
rect 6450 1950 6550 2050
rect 6650 1950 6750 2000
rect 6850 1950 6950 2000
rect 7050 1950 7150 2000
rect 7250 1950 7350 2000
rect 7450 1950 7550 2000
rect 7650 1950 7750 2000
rect 7850 1950 7950 2000
rect 8050 1950 8150 2000
rect 8250 1950 8350 2000
rect 8450 1950 8550 2000
rect 8650 1950 8750 2000
rect 8850 1950 8950 2000
rect 9050 1950 9150 2000
rect 9250 1950 9350 2050
rect 9454 2042 9478 2050
rect 9512 2042 9534 2076
rect 9454 2004 9534 2042
rect 9454 1970 9478 2004
rect 9512 1970 9534 2004
rect 9454 1950 9534 1970
rect 664 1932 9534 1950
rect 664 1898 688 1932
rect 722 1898 9478 1932
rect 9512 1898 9534 1932
rect 664 1860 9534 1898
rect 664 1826 688 1860
rect 722 1850 9478 1860
rect 722 1826 744 1850
rect 664 1788 744 1826
rect 664 1754 688 1788
rect 722 1754 744 1788
rect 664 1750 744 1754
rect 850 1750 950 1850
rect 1050 1750 1150 1850
rect 1250 1750 1350 1850
rect 1450 1750 1550 1850
rect 1650 1750 1750 1850
rect 1850 1750 1950 1850
rect 2050 1750 2150 1850
rect 2250 1750 2350 1850
rect 2450 1750 2550 1850
rect 2650 1750 2750 1850
rect 2850 1750 2950 1850
rect 3050 1750 3150 1850
rect 3250 1750 3350 1850
rect 3450 1750 3550 1850
rect 3650 1750 3750 1850
rect 3850 1750 3950 1850
rect 4050 1750 4150 1850
rect 4250 1750 4350 1850
rect 4450 1750 4550 1850
rect 4650 1750 4750 1850
rect 4850 1750 4950 1850
rect 5050 1750 5150 1850
rect 5250 1750 5350 1850
rect 5450 1750 5550 1850
rect 5650 1750 5750 1850
rect 5850 1750 5950 1850
rect 6050 1750 6150 1850
rect 6250 1750 6350 1850
rect 6450 1750 6550 1850
rect 6650 1750 6750 1850
rect 6850 1750 6950 1850
rect 7050 1750 7150 1850
rect 7250 1750 7350 1850
rect 7450 1750 7550 1850
rect 7650 1750 7750 1850
rect 7850 1750 7950 1850
rect 8050 1750 8150 1850
rect 8250 1750 8350 1850
rect 8450 1750 8550 1850
rect 8650 1750 8750 1850
rect 8850 1750 8950 1850
rect 9050 1750 9150 1850
rect 9250 1750 9350 1850
rect 9454 1826 9478 1850
rect 9512 1826 9534 1860
rect 9454 1788 9534 1826
rect 9454 1754 9478 1788
rect 9512 1754 9534 1788
rect 9454 1750 9534 1754
rect 664 1716 9534 1750
rect 664 1682 688 1716
rect 722 1682 9478 1716
rect 9512 1682 9534 1716
rect 664 1650 9534 1682
rect 664 1644 744 1650
rect 664 1610 688 1644
rect 722 1610 744 1644
rect 664 1572 744 1610
rect 664 1538 688 1572
rect 722 1550 744 1572
rect 850 1550 950 1650
rect 1050 1600 1150 1650
rect 1250 1600 1350 1650
rect 1450 1600 1550 1650
rect 1650 1600 1750 1650
rect 1850 1600 1950 1650
rect 2050 1600 2150 1650
rect 2250 1600 2350 1650
rect 2450 1600 2550 1650
rect 2650 1600 2750 1650
rect 2850 1600 2950 1650
rect 3050 1600 3150 1650
rect 3250 1600 3350 1650
rect 3450 1600 3550 1650
rect 3650 1550 3750 1650
rect 3850 1600 3950 1650
rect 4050 1600 4150 1650
rect 4250 1600 4350 1650
rect 4450 1600 4550 1650
rect 4650 1600 4750 1650
rect 4850 1600 4950 1650
rect 5050 1600 5150 1650
rect 5250 1600 5350 1650
rect 5450 1600 5550 1650
rect 5650 1600 5750 1650
rect 5850 1600 5950 1650
rect 6050 1600 6150 1650
rect 6250 1600 6350 1650
rect 6450 1550 6550 1650
rect 6650 1600 6750 1650
rect 6850 1600 6950 1650
rect 7050 1600 7150 1650
rect 7250 1600 7350 1650
rect 7450 1600 7550 1650
rect 7650 1600 7750 1650
rect 7850 1600 7950 1650
rect 8050 1600 8150 1650
rect 8250 1600 8350 1650
rect 8450 1600 8550 1650
rect 8650 1600 8750 1650
rect 8850 1600 8950 1650
rect 9050 1600 9150 1650
rect 9250 1550 9350 1650
rect 9454 1644 9534 1650
rect 9454 1610 9478 1644
rect 9512 1610 9534 1644
rect 9454 1572 9534 1610
rect 9454 1550 9478 1572
rect 722 1538 1000 1550
rect 664 1500 1000 1538
rect 664 1466 688 1500
rect 722 1466 1000 1500
rect 664 1450 1000 1466
rect 3600 1450 3800 1550
rect 6400 1450 6600 1550
rect 9200 1538 9478 1550
rect 9512 1538 9534 1572
rect 9200 1500 9534 1538
rect 9200 1466 9478 1500
rect 9512 1466 9534 1500
rect 9200 1450 9534 1466
rect 664 1428 744 1450
rect 664 1394 688 1428
rect 722 1394 744 1428
rect 664 1356 744 1394
rect 664 1322 688 1356
rect 722 1350 744 1356
rect 850 1350 950 1450
rect 722 1322 1000 1350
rect 664 1284 1000 1322
rect 664 1250 688 1284
rect 722 1250 1000 1284
rect 1122 1312 1202 1358
rect 1122 1278 1144 1312
rect 1178 1278 1202 1312
rect 664 1212 744 1250
rect 664 1178 688 1212
rect 722 1178 744 1212
rect 664 1150 744 1178
rect 850 1150 950 1250
rect 1122 1240 1202 1278
rect 1122 1206 1144 1240
rect 1178 1206 1202 1240
rect 1122 1168 1202 1206
rect 664 1140 1000 1150
rect 664 1106 688 1140
rect 722 1106 1000 1140
rect 664 1068 1000 1106
rect 664 1034 688 1068
rect 722 1050 1000 1068
rect 1122 1134 1144 1168
rect 1178 1134 1202 1168
rect 1122 1096 1202 1134
rect 1122 1062 1144 1096
rect 1178 1062 1202 1096
rect 722 1034 744 1050
rect 664 996 744 1034
rect 664 962 688 996
rect 722 962 744 996
rect 664 950 744 962
rect 850 950 950 1050
rect 1122 1024 1202 1062
rect 1122 990 1144 1024
rect 1178 990 1202 1024
rect 1122 952 1202 990
rect 664 924 1000 950
rect 664 890 688 924
rect 722 890 1000 924
rect 664 852 1000 890
rect 664 818 688 852
rect 722 850 1000 852
rect 1122 918 1144 952
rect 1178 918 1202 952
rect 1122 880 1202 918
rect 722 818 744 850
rect 664 780 744 818
rect 664 746 688 780
rect 722 746 744 780
rect 850 750 950 850
rect 1122 846 1144 880
rect 1178 846 1202 880
rect 1122 808 1202 846
rect 1122 774 1144 808
rect 1178 774 1202 808
rect 664 708 744 746
rect 800 650 1000 750
rect 1122 736 1202 774
rect 1122 702 1144 736
rect 1178 702 1202 736
rect 1122 664 1202 702
rect 50 550 150 650
rect 850 550 950 650
rect 1122 630 1144 664
rect 1178 630 1202 664
rect 1122 592 1202 630
rect 1122 558 1144 592
rect 1178 558 1202 592
rect 0 450 200 550
rect 800 450 1000 550
rect 1122 520 1202 558
rect 1122 486 1144 520
rect 1178 486 1202 520
rect 50 350 150 450
rect 250 350 350 400
rect 450 350 550 400
rect 650 350 750 400
rect 850 350 950 450
rect 1122 440 1202 486
rect 3398 1312 3478 1358
rect 3650 1350 3750 1450
rect 3398 1278 3420 1312
rect 3454 1278 3478 1312
rect 3398 1240 3478 1278
rect 3600 1250 3800 1350
rect 3922 1312 4000 1358
rect 3922 1278 3944 1312
rect 3978 1278 4000 1312
rect 3398 1206 3420 1240
rect 3454 1206 3478 1240
rect 3398 1168 3478 1206
rect 3398 1134 3420 1168
rect 3454 1134 3478 1168
rect 3650 1150 3750 1250
rect 3922 1240 4000 1278
rect 3922 1206 3944 1240
rect 3978 1206 4000 1240
rect 3922 1168 4000 1206
rect 3398 1096 3478 1134
rect 3398 1062 3420 1096
rect 3454 1062 3478 1096
rect 3398 1024 3478 1062
rect 3600 1050 3800 1150
rect 3922 1134 3944 1168
rect 3978 1134 4000 1168
rect 3922 1096 4000 1134
rect 3922 1062 3944 1096
rect 3978 1062 4000 1096
rect 3398 990 3420 1024
rect 3454 990 3478 1024
rect 3398 952 3478 990
rect 3398 918 3420 952
rect 3454 918 3478 952
rect 3650 950 3750 1050
rect 3922 1024 4000 1062
rect 3922 990 3944 1024
rect 3978 990 4000 1024
rect 3922 952 4000 990
rect 3398 880 3478 918
rect 3398 846 3420 880
rect 3454 846 3478 880
rect 3600 850 3800 950
rect 3922 918 3944 952
rect 3978 918 4000 952
rect 3922 880 4000 918
rect 3398 808 3478 846
rect 3398 774 3420 808
rect 3454 774 3478 808
rect 3398 736 3478 774
rect 3650 750 3750 850
rect 3922 846 3944 880
rect 3978 846 4000 880
rect 3922 808 4000 846
rect 3922 774 3944 808
rect 3978 774 4000 808
rect 3398 702 3420 736
rect 3454 702 3478 736
rect 3398 664 3478 702
rect 3398 630 3420 664
rect 3454 630 3478 664
rect 3600 650 3800 750
rect 3922 736 4000 774
rect 3922 702 3944 736
rect 3978 702 4000 736
rect 3922 664 4000 702
rect 3398 592 3478 630
rect 3398 558 3420 592
rect 3454 558 3478 592
rect 3398 520 3478 558
rect 3650 550 3750 650
rect 3922 630 3944 664
rect 3978 630 4000 664
rect 3922 592 4000 630
rect 3922 558 3944 592
rect 3978 558 4000 592
rect 3398 486 3420 520
rect 3454 486 3478 520
rect 3398 440 3478 486
rect 3600 450 3800 550
rect 3922 520 4000 558
rect 3922 486 3944 520
rect 3978 486 4000 520
rect 3650 350 3750 450
rect 3922 440 4000 486
rect 6198 1312 6278 1358
rect 6450 1350 6550 1450
rect 6198 1278 6220 1312
rect 6254 1278 6278 1312
rect 6198 1240 6278 1278
rect 6400 1250 6600 1350
rect 6722 1312 6802 1358
rect 6722 1278 6744 1312
rect 6778 1278 6802 1312
rect 6198 1206 6220 1240
rect 6254 1206 6278 1240
rect 6198 1168 6278 1206
rect 6198 1134 6220 1168
rect 6254 1134 6278 1168
rect 6450 1150 6550 1250
rect 6722 1240 6802 1278
rect 6722 1206 6744 1240
rect 6778 1206 6802 1240
rect 6722 1168 6802 1206
rect 6198 1096 6278 1134
rect 6198 1062 6220 1096
rect 6254 1062 6278 1096
rect 6198 1024 6278 1062
rect 6400 1050 6600 1150
rect 6722 1134 6744 1168
rect 6778 1134 6802 1168
rect 6722 1096 6802 1134
rect 6722 1062 6744 1096
rect 6778 1062 6802 1096
rect 6198 990 6220 1024
rect 6254 990 6278 1024
rect 6198 952 6278 990
rect 6198 918 6220 952
rect 6254 918 6278 952
rect 6450 950 6550 1050
rect 6722 1024 6802 1062
rect 6722 990 6744 1024
rect 6778 990 6802 1024
rect 6722 952 6802 990
rect 6198 880 6278 918
rect 6198 846 6220 880
rect 6254 846 6278 880
rect 6400 850 6600 950
rect 6722 918 6744 952
rect 6778 918 6802 952
rect 6722 880 6802 918
rect 6198 808 6278 846
rect 6198 774 6220 808
rect 6254 774 6278 808
rect 6198 736 6278 774
rect 6450 750 6550 850
rect 6722 846 6744 880
rect 6778 846 6802 880
rect 6722 808 6802 846
rect 6722 774 6744 808
rect 6778 774 6802 808
rect 6198 702 6220 736
rect 6254 702 6278 736
rect 6198 664 6278 702
rect 6198 630 6220 664
rect 6254 630 6278 664
rect 6400 650 6600 750
rect 6722 736 6802 774
rect 6722 702 6744 736
rect 6778 702 6802 736
rect 6722 664 6802 702
rect 6198 592 6278 630
rect 6198 558 6220 592
rect 6254 558 6278 592
rect 6198 520 6278 558
rect 6450 550 6550 650
rect 6722 630 6744 664
rect 6778 630 6802 664
rect 6722 592 6802 630
rect 6722 558 6744 592
rect 6778 558 6802 592
rect 6198 486 6220 520
rect 6254 486 6278 520
rect 6198 440 6278 486
rect 6400 450 6600 550
rect 6722 520 6802 558
rect 6722 486 6744 520
rect 6778 486 6802 520
rect 6450 350 6550 450
rect 6722 440 6802 486
rect 8996 1312 9078 1358
rect 9250 1350 9350 1450
rect 9454 1428 9534 1450
rect 9454 1394 9478 1428
rect 9512 1394 9534 1428
rect 9454 1356 9534 1394
rect 9454 1350 9478 1356
rect 8996 1278 9020 1312
rect 9054 1278 9078 1312
rect 8996 1240 9078 1278
rect 9200 1322 9478 1350
rect 9512 1322 9534 1356
rect 9200 1284 9534 1322
rect 9200 1250 9478 1284
rect 9512 1250 9534 1284
rect 8996 1206 9020 1240
rect 9054 1206 9078 1240
rect 8996 1168 9078 1206
rect 8996 1134 9020 1168
rect 9054 1134 9078 1168
rect 9250 1150 9350 1250
rect 9454 1212 9534 1250
rect 9454 1178 9478 1212
rect 9512 1178 9534 1212
rect 9454 1150 9534 1178
rect 8996 1096 9078 1134
rect 8996 1062 9020 1096
rect 9054 1062 9078 1096
rect 8996 1024 9078 1062
rect 9200 1140 9534 1150
rect 9200 1106 9478 1140
rect 9512 1106 9534 1140
rect 9200 1068 9534 1106
rect 9200 1050 9478 1068
rect 8996 990 9020 1024
rect 9054 990 9078 1024
rect 8996 952 9078 990
rect 8996 918 9020 952
rect 9054 918 9078 952
rect 9250 950 9350 1050
rect 9454 1034 9478 1050
rect 9512 1034 9534 1068
rect 9454 996 9534 1034
rect 9454 962 9478 996
rect 9512 962 9534 996
rect 9454 950 9534 962
rect 8996 880 9078 918
rect 8996 846 9020 880
rect 9054 846 9078 880
rect 9200 924 9534 950
rect 9200 890 9478 924
rect 9512 890 9534 924
rect 9200 852 9534 890
rect 9200 850 9478 852
rect 8996 808 9078 846
rect 8996 774 9020 808
rect 9054 774 9078 808
rect 8996 736 9078 774
rect 9250 750 9350 850
rect 9454 818 9478 850
rect 9512 818 9534 852
rect 9454 780 9534 818
rect 8996 702 9020 736
rect 9054 702 9078 736
rect 8996 664 9078 702
rect 8996 630 9020 664
rect 9054 630 9078 664
rect 9200 650 9400 750
rect 9454 746 9478 780
rect 9512 746 9534 780
rect 9454 708 9534 746
rect 9864 2618 9888 2652
rect 9922 2618 9944 2652
rect 10000 2650 10200 2750
rect 9864 2580 9944 2618
rect 9864 2546 9888 2580
rect 9922 2550 9944 2580
rect 10050 2550 10150 2650
rect 9922 2546 10200 2550
rect 9864 2508 10200 2546
rect 9864 2474 9888 2508
rect 9922 2474 10200 2508
rect 9864 2450 10200 2474
rect 9864 2436 9944 2450
rect 9864 2402 9888 2436
rect 9922 2402 9944 2436
rect 9864 2364 9944 2402
rect 9864 2330 9888 2364
rect 9922 2350 9944 2364
rect 10050 2350 10150 2450
rect 9922 2330 10200 2350
rect 9864 2292 10200 2330
rect 9864 2258 9888 2292
rect 9922 2258 10200 2292
rect 9864 2250 10200 2258
rect 9864 2220 9944 2250
rect 9864 2186 9888 2220
rect 9922 2186 9944 2220
rect 9864 2150 9944 2186
rect 10050 2150 10150 2250
rect 9864 2148 10200 2150
rect 9864 2114 9888 2148
rect 9922 2114 10200 2148
rect 9864 2076 10200 2114
rect 9864 2042 9888 2076
rect 9922 2050 10200 2076
rect 9922 2042 9944 2050
rect 9864 2004 9944 2042
rect 9864 1970 9888 2004
rect 9922 1970 9944 2004
rect 9864 1950 9944 1970
rect 10050 1950 10150 2050
rect 9864 1932 10200 1950
rect 9864 1898 9888 1932
rect 9922 1898 10200 1932
rect 9864 1860 10200 1898
rect 9864 1826 9888 1860
rect 9922 1850 10200 1860
rect 9922 1826 9944 1850
rect 9864 1788 9944 1826
rect 9864 1754 9888 1788
rect 9922 1754 9944 1788
rect 9864 1750 9944 1754
rect 10050 1750 10150 1850
rect 9864 1716 10200 1750
rect 9864 1682 9888 1716
rect 9922 1682 10200 1716
rect 9864 1650 10200 1682
rect 9864 1644 9944 1650
rect 9864 1610 9888 1644
rect 9922 1610 9944 1644
rect 9864 1572 9944 1610
rect 9864 1538 9888 1572
rect 9922 1550 9944 1572
rect 10050 1550 10150 1650
rect 9922 1538 10200 1550
rect 9864 1500 10200 1538
rect 9864 1466 9888 1500
rect 9922 1466 10200 1500
rect 9864 1450 10200 1466
rect 9864 1428 9944 1450
rect 9864 1394 9888 1428
rect 9922 1394 9944 1428
rect 9864 1356 9944 1394
rect 9864 1322 9888 1356
rect 9922 1350 9944 1356
rect 10050 1350 10150 1450
rect 9922 1322 10200 1350
rect 9864 1284 10200 1322
rect 9864 1250 9888 1284
rect 9922 1250 10200 1284
rect 9864 1212 9944 1250
rect 9864 1178 9888 1212
rect 9922 1178 9944 1212
rect 9864 1150 9944 1178
rect 10050 1150 10150 1250
rect 9864 1140 10200 1150
rect 9864 1106 9888 1140
rect 9922 1106 10200 1140
rect 9864 1068 10200 1106
rect 9864 1034 9888 1068
rect 9922 1050 10200 1068
rect 9922 1034 9944 1050
rect 9864 996 9944 1034
rect 9864 962 9888 996
rect 9922 962 9944 996
rect 9864 950 9944 962
rect 10050 950 10150 1050
rect 9864 924 10200 950
rect 9864 890 9888 924
rect 9922 890 10200 924
rect 9864 852 10200 890
rect 9864 818 9888 852
rect 9922 850 10200 852
rect 9922 818 9944 850
rect 9864 780 9944 818
rect 9864 746 9888 780
rect 9922 746 9944 780
rect 10050 750 10150 850
rect 9864 708 9944 746
rect 10000 650 10200 750
rect 8996 592 9078 630
rect 8996 558 9020 592
rect 9054 558 9078 592
rect 8996 520 9078 558
rect 9250 550 9350 650
rect 10050 550 10150 650
rect 8996 486 9020 520
rect 9054 486 9078 520
rect 8996 440 9078 486
rect 9200 450 9400 550
rect 10000 450 10200 550
rect 9250 350 9350 450
rect 9450 350 9550 400
rect 9650 350 9750 400
rect 9850 350 9950 400
rect 10050 350 10150 450
rect 0 250 1000 350
rect 3600 250 3800 350
rect 6400 250 6600 350
rect 9200 250 10200 350
rect 50 150 150 250
rect 250 150 350 250
rect 450 150 550 250
rect 650 150 750 250
rect 850 150 950 250
rect 1050 150 1150 200
rect 1250 150 1350 200
rect 1450 150 1550 200
rect 1650 150 1750 200
rect 1850 150 1950 200
rect 2050 150 2150 200
rect 2250 150 2350 200
rect 2450 150 2550 200
rect 2650 150 2750 200
rect 2850 150 2950 200
rect 3050 150 3150 200
rect 3250 150 3350 200
rect 3450 150 3550 200
rect 3650 150 3750 250
rect 3850 150 3950 200
rect 4050 150 4150 200
rect 4250 150 4350 200
rect 4450 150 4550 200
rect 4650 150 4750 200
rect 4850 150 4950 200
rect 5050 150 5150 200
rect 5250 150 5350 200
rect 5450 150 5550 200
rect 5650 150 5750 200
rect 5850 150 5950 200
rect 6050 150 6150 200
rect 6250 150 6350 200
rect 6450 150 6550 250
rect 6650 150 6750 200
rect 6850 150 6950 200
rect 7050 150 7150 200
rect 7250 150 7350 200
rect 7450 150 7550 200
rect 7650 150 7750 200
rect 7850 150 7950 200
rect 8050 150 8150 200
rect 8250 150 8350 200
rect 8450 150 8550 200
rect 8650 150 8750 200
rect 8850 150 8950 200
rect 9050 150 9150 200
rect 9250 150 9350 250
rect 9450 150 9550 250
rect 9650 150 9750 250
rect 9850 150 9950 250
rect 10050 150 10150 250
rect 0 50 10200 150
rect 50 0 150 50
rect 250 0 350 50
rect 450 0 550 50
rect 650 0 750 50
rect 850 0 950 50
rect 1050 0 1150 50
rect 1250 0 1350 50
rect 1450 0 1550 50
rect 1650 0 1750 50
rect 1850 0 1950 50
rect 2050 0 2150 50
rect 2250 0 2350 50
rect 2450 0 2550 50
rect 2650 0 2750 50
rect 2850 0 2950 50
rect 3050 0 3150 50
rect 3250 0 3350 50
rect 3450 0 3550 50
rect 3650 0 3750 50
rect 3850 0 3950 50
rect 4050 0 4150 50
rect 4250 0 4350 50
rect 4450 0 4550 50
rect 4650 0 4750 50
rect 4850 0 4950 50
rect 5050 0 5150 50
rect 5250 0 5350 50
rect 5450 0 5550 50
rect 5650 0 5750 50
rect 5850 0 5950 50
rect 6050 0 6150 50
rect 6250 0 6350 50
rect 6450 0 6550 50
rect 6650 0 6750 50
rect 6850 0 6950 50
rect 7050 0 7150 50
rect 7250 0 7350 50
rect 7450 0 7550 50
rect 7650 0 7750 50
rect 7850 0 7950 50
rect 8050 0 8150 50
rect 8250 0 8350 50
rect 8450 0 8550 50
rect 8650 0 8750 50
rect 8850 0 8950 50
rect 9050 0 9150 50
rect 9250 0 9350 50
rect 9450 0 9550 50
rect 9650 0 9750 50
rect 9850 0 9950 50
rect 10050 0 10150 50
<< metal2 >>
rect 50 3550 150 3600
rect 250 3550 350 3600
rect 450 3550 550 3600
rect 650 3550 750 3600
rect 850 3550 950 3600
rect 1050 3550 1150 3600
rect 1250 3550 1350 3600
rect 1450 3550 1550 3600
rect 1650 3550 1750 3600
rect 1850 3550 1950 3600
rect 2050 3550 2150 3600
rect 2250 3550 2350 3600
rect 2450 3550 2550 3600
rect 2650 3550 2750 3600
rect 2850 3550 2950 3600
rect 3050 3550 3150 3600
rect 3250 3550 3350 3600
rect 3450 3550 3550 3600
rect 3650 3550 3750 3600
rect 3850 3550 3950 3600
rect 4050 3550 4150 3600
rect 4250 3550 4350 3600
rect 4450 3550 4550 3600
rect 4650 3550 4750 3600
rect 4850 3550 4950 3600
rect 5050 3550 5150 3600
rect 5250 3550 5350 3600
rect 5450 3550 5550 3600
rect 5650 3550 5750 3600
rect 5850 3550 5950 3600
rect 6050 3550 6150 3600
rect 6250 3550 6350 3600
rect 6450 3550 6550 3600
rect 6650 3550 6750 3600
rect 6850 3550 6950 3600
rect 7050 3550 7150 3600
rect 7250 3550 7350 3600
rect 7450 3550 7550 3600
rect 7650 3550 7750 3600
rect 7850 3550 7950 3600
rect 8050 3550 8150 3600
rect 8250 3550 8350 3600
rect 8450 3550 8550 3600
rect 8650 3550 8750 3600
rect 8850 3550 8950 3600
rect 9050 3550 9150 3600
rect 9250 3550 9350 3600
rect 9450 3550 9550 3600
rect 9650 3550 9750 3600
rect 9850 3550 9950 3600
rect 10050 3550 10150 3600
rect 0 3450 10200 3550
rect 50 3350 150 3450
rect 250 3350 350 3450
rect 450 3350 550 3450
rect 650 3350 750 3450
rect 850 3350 950 3450
rect 1050 3400 1150 3450
rect 1250 3400 1350 3450
rect 1450 3400 1550 3450
rect 1650 3400 1750 3450
rect 1850 3400 1950 3450
rect 2050 3400 2150 3450
rect 2250 3400 2350 3450
rect 2450 3400 2550 3450
rect 2650 3400 2750 3450
rect 2850 3400 2950 3450
rect 3050 3400 3150 3450
rect 3250 3400 3350 3450
rect 3450 3400 3550 3450
rect 3650 3350 3750 3450
rect 3850 3400 3950 3450
rect 4050 3400 4150 3450
rect 4250 3400 4350 3450
rect 4450 3400 4550 3450
rect 4650 3400 4750 3450
rect 4850 3400 4950 3450
rect 5050 3400 5150 3450
rect 5250 3400 5350 3450
rect 5450 3400 5550 3450
rect 5650 3400 5750 3450
rect 5850 3400 5950 3450
rect 6050 3400 6150 3450
rect 6250 3400 6350 3450
rect 6450 3350 6550 3450
rect 6650 3400 6750 3450
rect 6850 3400 6950 3450
rect 7050 3400 7150 3450
rect 7250 3400 7350 3450
rect 7450 3400 7550 3450
rect 7650 3400 7750 3450
rect 7850 3400 7950 3450
rect 8050 3400 8150 3450
rect 8250 3400 8350 3450
rect 8450 3400 8550 3450
rect 8650 3400 8750 3450
rect 8850 3400 8950 3450
rect 9050 3400 9150 3450
rect 9250 3350 9350 3450
rect 9450 3350 9550 3450
rect 9650 3350 9750 3450
rect 9850 3350 9950 3450
rect 10050 3350 10150 3450
rect 0 3250 1000 3350
rect 3600 3250 3800 3350
rect 6400 3250 6600 3350
rect 9200 3250 10200 3350
rect 50 3150 150 3250
rect 250 3150 350 3250
rect 450 3150 550 3250
rect 650 3150 750 3250
rect 850 3150 950 3250
rect 1122 3150 1202 3158
rect 0 3050 1202 3150
rect 50 2950 150 3050
rect 250 3000 350 3050
rect 450 3000 550 3050
rect 650 3000 750 3050
rect 850 2950 950 3050
rect 1122 2950 1202 3050
rect 0 2850 200 2950
rect 800 2850 1202 2950
rect 50 2750 150 2850
rect 0 2650 200 2750
rect 50 2550 150 2650
rect 0 2450 200 2550
rect 50 2350 150 2450
rect 450 2400 550 2800
rect 850 2750 950 2850
rect 1122 2750 1202 2850
rect 800 2650 1202 2750
rect 850 2550 950 2650
rect 1122 2550 1202 2650
rect 800 2450 1202 2550
rect 850 2350 950 2450
rect 1122 2350 1202 2450
rect 0 2250 200 2350
rect 800 2250 1202 2350
rect 50 2150 150 2250
rect 850 2150 950 2250
rect 1122 2240 1202 2250
rect 3398 3150 3478 3158
rect 3650 3150 3750 3250
rect 3922 3150 4000 3158
rect 3398 3050 4000 3150
rect 3398 2950 3478 3050
rect 3650 2950 3750 3050
rect 3922 2950 4000 3050
rect 3398 2850 4000 2950
rect 3398 2750 3478 2850
rect 3650 2750 3750 2850
rect 3922 2750 4000 2850
rect 3398 2650 4000 2750
rect 3398 2550 3478 2650
rect 3650 2550 3750 2650
rect 3922 2550 4000 2650
rect 3398 2450 4000 2550
rect 3398 2350 3478 2450
rect 3650 2350 3750 2450
rect 3922 2350 4000 2450
rect 3398 2250 4000 2350
rect 6198 3150 6278 3158
rect 6450 3150 6550 3250
rect 6722 3150 6802 3158
rect 6198 3050 6802 3150
rect 6198 2950 6278 3050
rect 6450 2950 6550 3050
rect 6722 2950 6802 3050
rect 6198 2850 6802 2950
rect 6198 2750 6278 2850
rect 6450 2750 6550 2850
rect 6722 2750 6802 2850
rect 6198 2650 6802 2750
rect 6198 2550 6278 2650
rect 6450 2550 6550 2650
rect 6722 2550 6802 2650
rect 6198 2450 6802 2550
rect 6198 2350 6278 2450
rect 6450 2350 6550 2450
rect 6722 2350 6802 2450
rect 3398 2240 3478 2250
rect 3650 2150 3750 2250
rect 3922 2240 4000 2250
rect 0 2050 200 2150
rect 800 2050 1000 2150
rect 3600 2050 3800 2150
rect 50 1950 150 2050
rect 850 1950 950 2050
rect 1050 1950 1150 2000
rect 1250 1950 1350 2000
rect 1450 1950 1550 2000
rect 1650 1950 1750 2000
rect 1850 1950 1950 2000
rect 2050 1950 2150 2000
rect 2250 1950 2350 2000
rect 2450 1950 2550 2000
rect 2650 1950 2750 2000
rect 2850 1950 2950 2000
rect 3050 1950 3150 2000
rect 3250 1950 3350 2000
rect 3450 1950 3550 2000
rect 3650 1950 3750 2050
rect 3850 1950 3950 2000
rect 4050 1950 4150 2000
rect 4250 1950 4350 2300
rect 4450 1950 4550 2300
rect 4650 1950 4750 2300
rect 4850 1950 4950 2300
rect 5050 1950 5150 2300
rect 5250 1950 5350 2300
rect 5450 1950 5550 2300
rect 5650 1950 5750 2300
rect 5850 1950 5950 2300
rect 6198 2250 6802 2350
rect 6198 2240 6278 2250
rect 6450 2150 6550 2250
rect 6722 2240 6802 2250
rect 8996 3150 9078 3158
rect 9250 3150 9350 3250
rect 9450 3150 9550 3250
rect 9650 3150 9750 3250
rect 9850 3150 9950 3250
rect 10050 3150 10150 3250
rect 8996 3050 10200 3150
rect 8996 2950 9078 3050
rect 9250 2950 9350 3050
rect 9450 3000 9550 3050
rect 9650 3000 9750 3050
rect 9850 3000 9950 3050
rect 10050 2950 10150 3050
rect 8996 2850 9400 2950
rect 10000 2850 10200 2950
rect 8996 2750 9078 2850
rect 9250 2750 9350 2850
rect 8996 2650 9400 2750
rect 8996 2550 9078 2650
rect 9250 2550 9350 2650
rect 8996 2450 9400 2550
rect 8996 2350 9078 2450
rect 9250 2350 9350 2450
rect 9650 2400 9750 2800
rect 10050 2750 10150 2850
rect 10000 2650 10200 2750
rect 10050 2550 10150 2650
rect 10000 2450 10200 2550
rect 10050 2350 10150 2450
rect 8996 2250 9400 2350
rect 10000 2250 10200 2350
rect 8996 2240 9078 2250
rect 9250 2150 9350 2250
rect 10050 2150 10150 2250
rect 6400 2050 6600 2150
rect 9200 2050 9400 2150
rect 10000 2050 10200 2150
rect 6050 1950 6150 2000
rect 6250 1950 6350 2000
rect 6450 1950 6550 2050
rect 6650 1950 6750 2000
rect 6850 1950 6950 2000
rect 7050 1950 7150 2000
rect 7250 1950 7350 2000
rect 7450 1950 7550 2000
rect 7650 1950 7750 2000
rect 7850 1950 7950 2000
rect 8050 1950 8150 2000
rect 8250 1950 8350 2000
rect 8450 1950 8550 2000
rect 8650 1950 8750 2000
rect 8850 1950 8950 2000
rect 9050 1950 9150 2000
rect 9250 1950 9350 2050
rect 10050 1950 10150 2050
rect 0 1850 200 1950
rect 800 1850 9400 1950
rect 10000 1850 10200 1950
rect 50 1750 150 1850
rect 850 1750 950 1850
rect 1050 1750 1150 1850
rect 1250 1750 1350 1850
rect 1450 1750 1550 1850
rect 1650 1750 1750 1850
rect 1850 1750 1950 1850
rect 2050 1750 2150 1850
rect 2250 1750 2350 1850
rect 2450 1750 2550 1850
rect 2650 1750 2750 1850
rect 2850 1750 2950 1850
rect 3050 1750 3150 1850
rect 3250 1750 3350 1850
rect 3450 1750 3550 1850
rect 3650 1750 3750 1850
rect 3850 1750 3950 1850
rect 4050 1750 4150 1850
rect 4250 1750 4350 1850
rect 4450 1750 4550 1850
rect 4650 1750 4750 1850
rect 4850 1750 4950 1850
rect 5050 1750 5150 1850
rect 5250 1750 5350 1850
rect 5450 1750 5550 1850
rect 5650 1750 5750 1850
rect 5850 1750 5950 1850
rect 6050 1750 6150 1850
rect 6250 1750 6350 1850
rect 6450 1750 6550 1850
rect 6650 1750 6750 1850
rect 6850 1750 6950 1850
rect 7050 1750 7150 1850
rect 7250 1750 7350 1850
rect 7450 1750 7550 1850
rect 7650 1750 7750 1850
rect 7850 1750 7950 1850
rect 8050 1750 8150 1850
rect 8250 1750 8350 1850
rect 8450 1750 8550 1850
rect 8650 1750 8750 1850
rect 8850 1750 8950 1850
rect 9050 1750 9150 1850
rect 9250 1750 9350 1850
rect 10050 1750 10150 1850
rect 0 1650 200 1750
rect 800 1650 9400 1750
rect 10000 1650 10200 1750
rect 50 1550 150 1650
rect 850 1550 950 1650
rect 1050 1600 1150 1650
rect 1250 1600 1350 1650
rect 1450 1600 1550 1650
rect 1650 1600 1750 1650
rect 1850 1600 1950 1650
rect 2050 1600 2150 1650
rect 2250 1600 2350 1650
rect 2450 1600 2550 1650
rect 2650 1600 2750 1650
rect 2850 1600 2950 1650
rect 3050 1600 3150 1650
rect 3250 1600 3350 1650
rect 3450 1600 3550 1650
rect 3650 1550 3750 1650
rect 3850 1600 3950 1650
rect 4050 1600 4150 1650
rect 0 1450 200 1550
rect 800 1450 1000 1550
rect 3600 1450 3800 1550
rect 50 1350 150 1450
rect 850 1350 950 1450
rect 1122 1350 1202 1358
rect 0 1250 200 1350
rect 800 1250 1202 1350
rect 50 1150 150 1250
rect 850 1150 950 1250
rect 1122 1150 1202 1250
rect 0 1050 200 1150
rect 800 1050 1202 1150
rect 50 950 150 1050
rect 850 950 950 1050
rect 1122 950 1202 1050
rect 0 850 200 950
rect 800 850 1202 950
rect 50 750 150 850
rect 850 750 950 850
rect 1122 750 1202 850
rect 0 650 200 750
rect 800 650 1202 750
rect 50 550 150 650
rect 850 550 950 650
rect 1122 550 1202 650
rect 0 450 200 550
rect 800 450 1202 550
rect 50 350 150 450
rect 250 350 350 400
rect 450 350 550 400
rect 650 350 750 400
rect 850 350 950 450
rect 1122 440 1202 450
rect 3398 1350 3478 1358
rect 3650 1350 3750 1450
rect 3922 1350 4000 1358
rect 3398 1250 4000 1350
rect 3398 1150 3478 1250
rect 3650 1150 3750 1250
rect 3922 1150 4000 1250
rect 4250 1200 4350 1650
rect 4450 1200 4550 1650
rect 4650 1200 4750 1650
rect 4850 1200 4950 1650
rect 5050 1200 5150 1650
rect 5250 1200 5350 1650
rect 5450 1200 5550 1650
rect 5650 1200 5750 1650
rect 5850 1200 5950 1650
rect 6050 1600 6150 1650
rect 6250 1600 6350 1650
rect 6450 1550 6550 1650
rect 6650 1600 6750 1650
rect 6850 1600 6950 1650
rect 7050 1600 7150 1650
rect 7250 1600 7350 1650
rect 7450 1600 7550 1650
rect 7650 1600 7750 1650
rect 7850 1600 7950 1650
rect 8050 1600 8150 1650
rect 8250 1600 8350 1650
rect 8450 1600 8550 1650
rect 8650 1600 8750 1650
rect 8850 1600 8950 1650
rect 9050 1600 9150 1650
rect 9250 1550 9350 1650
rect 10050 1550 10150 1650
rect 6400 1450 6600 1550
rect 9200 1450 9400 1550
rect 10000 1450 10200 1550
rect 6198 1350 6278 1358
rect 6450 1350 6550 1450
rect 6722 1350 6802 1358
rect 6198 1250 6802 1350
rect 3398 1050 4000 1150
rect 3398 950 3478 1050
rect 3650 950 3750 1050
rect 3922 950 4000 1050
rect 3398 850 4000 950
rect 3398 750 3478 850
rect 3650 750 3750 850
rect 3922 750 4000 850
rect 3398 650 4000 750
rect 3398 550 3478 650
rect 3650 550 3750 650
rect 3922 550 4000 650
rect 3398 450 4000 550
rect 3398 440 3478 450
rect 3650 350 3750 450
rect 3922 440 4000 450
rect 6198 1150 6278 1250
rect 6450 1150 6550 1250
rect 6722 1150 6802 1250
rect 6198 1050 6802 1150
rect 6198 950 6278 1050
rect 6450 950 6550 1050
rect 6722 950 6802 1050
rect 6198 850 6802 950
rect 6198 750 6278 850
rect 6450 750 6550 850
rect 6722 750 6802 850
rect 6198 650 6802 750
rect 6198 550 6278 650
rect 6450 550 6550 650
rect 6722 550 6802 650
rect 6198 450 6802 550
rect 6198 440 6278 450
rect 6450 350 6550 450
rect 6722 440 6802 450
rect 8996 1350 9078 1358
rect 9250 1350 9350 1450
rect 10050 1350 10150 1450
rect 8996 1250 9400 1350
rect 10000 1250 10200 1350
rect 8996 1150 9078 1250
rect 9250 1150 9350 1250
rect 10050 1150 10150 1250
rect 8996 1050 9400 1150
rect 10000 1050 10200 1150
rect 8996 950 9078 1050
rect 9250 950 9350 1050
rect 10050 950 10150 1050
rect 8996 850 9400 950
rect 10000 850 10200 950
rect 8996 750 9078 850
rect 9250 750 9350 850
rect 10050 750 10150 850
rect 8996 650 9400 750
rect 10000 650 10200 750
rect 8996 550 9078 650
rect 9250 550 9350 650
rect 10050 550 10150 650
rect 8996 450 9400 550
rect 10000 450 10200 550
rect 8996 440 9078 450
rect 9250 350 9350 450
rect 9450 350 9550 400
rect 9650 350 9750 400
rect 9850 350 9950 400
rect 10050 350 10150 450
rect 0 250 1000 350
rect 3600 250 3800 350
rect 6400 250 6600 350
rect 9200 250 10200 350
rect 50 150 150 250
rect 250 150 350 250
rect 450 150 550 250
rect 650 150 750 250
rect 850 150 950 250
rect 1050 150 1150 200
rect 1250 150 1350 200
rect 1450 150 1550 200
rect 1650 150 1750 200
rect 1850 150 1950 200
rect 2050 150 2150 200
rect 2250 150 2350 200
rect 2450 150 2550 200
rect 2650 150 2750 200
rect 2850 150 2950 200
rect 3050 150 3150 200
rect 3250 150 3350 200
rect 3450 150 3550 200
rect 3650 150 3750 250
rect 3850 150 3950 200
rect 4050 150 4150 200
rect 4250 150 4350 200
rect 4450 150 4550 200
rect 4650 150 4750 200
rect 4850 150 4950 200
rect 5050 150 5150 200
rect 5250 150 5350 200
rect 5450 150 5550 200
rect 5650 150 5750 200
rect 5850 150 5950 200
rect 6050 150 6150 200
rect 6250 150 6350 200
rect 6450 150 6550 250
rect 6650 150 6750 200
rect 6850 150 6950 200
rect 7050 150 7150 200
rect 7250 150 7350 200
rect 7450 150 7550 200
rect 7650 150 7750 200
rect 7850 150 7950 200
rect 8050 150 8150 200
rect 8250 150 8350 200
rect 8450 150 8550 200
rect 8650 150 8750 200
rect 8850 150 8950 200
rect 9050 150 9150 200
rect 9250 150 9350 250
rect 9450 150 9550 250
rect 9650 150 9750 250
rect 9850 150 9950 250
rect 10050 150 10150 250
rect 0 50 10200 150
rect 50 0 150 50
rect 250 0 350 50
rect 450 0 550 50
rect 650 0 750 50
rect 850 0 950 50
rect 1050 0 1150 50
rect 1250 0 1350 50
rect 1450 0 1550 50
rect 1650 0 1750 50
rect 1850 0 1950 50
rect 2050 0 2150 50
rect 2250 0 2350 50
rect 2450 0 2550 50
rect 2650 0 2750 50
rect 2850 0 2950 50
rect 3050 0 3150 50
rect 3250 0 3350 50
rect 3450 0 3550 50
rect 3650 0 3750 50
rect 3850 0 3950 50
rect 4050 0 4150 50
rect 4250 0 4350 50
rect 4450 0 4550 50
rect 4650 0 4750 50
rect 4850 0 4950 50
rect 5050 0 5150 50
rect 5250 0 5350 50
rect 5450 0 5550 50
rect 5650 0 5750 50
rect 5850 0 5950 50
rect 6050 0 6150 50
rect 6250 0 6350 50
rect 6450 0 6550 50
rect 6650 0 6750 50
rect 6850 0 6950 50
rect 7050 0 7150 50
rect 7250 0 7350 50
rect 7450 0 7550 50
rect 7650 0 7750 50
rect 7850 0 7950 50
rect 8050 0 8150 50
rect 8250 0 8350 50
rect 8450 0 8550 50
rect 8650 0 8750 50
rect 8850 0 8950 50
rect 9050 0 9150 50
rect 9250 0 9350 50
rect 9450 0 9550 50
rect 9650 0 9750 50
rect 9850 0 9950 50
rect 10050 0 10150 50
<< metal3 >>
rect 2250 2650 2350 2750
rect 4050 2740 4150 2750
rect 3060 2660 4150 2740
rect 2260 950 2340 2650
rect 3060 2350 3140 2660
rect 4050 2650 4150 2660
rect 6050 2740 6150 2750
rect 6050 2660 7140 2740
rect 6050 2650 6150 2660
rect 7060 2350 7140 2660
rect 7850 2650 7950 2750
rect 3050 2250 3150 2350
rect 7050 2250 7150 2350
rect 3050 1250 3150 1350
rect 7050 1340 7150 1350
rect 3260 1260 7150 1340
rect 3060 1150 3140 1250
rect 3050 1050 3150 1150
rect 3260 950 3340 1260
rect 7050 1250 7150 1260
rect 7860 950 7940 2650
rect 450 940 550 950
rect 1250 940 1350 950
rect 450 860 1350 940
rect 450 850 550 860
rect 1250 850 1350 860
rect 2250 850 2350 950
rect 3250 850 3350 950
rect 4050 850 4150 950
rect 6050 850 6150 950
rect 6650 940 6750 950
rect 6850 940 6950 950
rect 6650 860 6950 940
rect 6650 850 6750 860
rect 6850 850 6950 860
rect 7850 850 7950 950
rect 8850 940 8950 950
rect 9650 940 9750 950
rect 8850 860 9750 940
rect 8850 850 8950 860
rect 9650 850 9750 860
rect 4060 740 4140 850
rect 3460 660 4140 740
rect 6060 740 6140 850
rect 6060 660 6740 740
rect 3050 540 3150 550
rect 3460 540 3540 660
rect 3050 460 3540 540
rect 6660 540 6740 660
rect 7050 540 7150 550
rect 6660 460 7150 540
rect 3050 450 3150 460
rect 7050 450 7150 460
<< metal4 >>
rect 3060 1060 6740 1140
rect 6660 860 6740 1060
use via_M1_M2_1_a  NoName_203 ~/A2G/MAGIC/magic_layout/skywater130_microtemplates_dense
timestamp 1647525606
transform 1 0 1162 0 1 2700
box -32 -32 32 32
use via_M1_M2_1_b  NoName_204 ~/A2G/MAGIC/magic_layout/skywater130_microtemplates_dense
timestamp 1647525606
transform 1 0 1162 0 1 2828
box -32 -32 32 32
use via_M1_M2_1_c  NoName_205 ~/A2G/MAGIC/magic_layout/skywater130_microtemplates_dense
timestamp 1647525606
transform 1 0 1162 0 1 2572
box -32 -32 32 32
use via_M1_M2_1_d  NoName_206 ~/A2G/MAGIC/magic_layout/skywater130_microtemplates_dense
timestamp 1647525606
transform 1 0 1162 0 1 2956
box -32 -32 32 32
use via_M1_M2_1_e  NoName_207 ~/A2G/MAGIC/magic_layout/skywater130_microtemplates_dense
timestamp 1647525606
transform 1 0 1162 0 1 2444
box -32 -32 32 32
use via_M1_M2_1_f  NoName_208 ~/A2G/MAGIC/magic_layout/skywater130_microtemplates_dense
timestamp 1647525606
transform 1 0 1162 0 1 3084
box -32 -32 32 32
use via_M1_M2_1_g  NoName_209 ~/A2G/MAGIC/magic_layout/skywater130_microtemplates_dense
timestamp 1647525606
transform 1 0 1162 0 1 2316
box -32 -32 32 32
use via_M1_M2_1_h  NoName_210 ~/A2G/MAGIC/magic_layout/skywater130_microtemplates_dense
timestamp 1647525606
transform 1 0 3438 0 1 2700
box -32 -32 32 32
use via_M1_M2_1_i  NoName_211 ~/A2G/MAGIC/magic_layout/skywater130_microtemplates_dense
timestamp 1647525606
transform 1 0 3438 0 1 2828
box -32 -32 32 32
use via_M1_M2_1_j  NoName_212 ~/A2G/MAGIC/magic_layout/skywater130_microtemplates_dense
timestamp 1647525606
transform 1 0 3438 0 1 2572
box -32 -32 32 32
use via_M1_M2_1_k  NoName_213 ~/A2G/MAGIC/magic_layout/skywater130_microtemplates_dense
timestamp 1647525606
transform 1 0 3438 0 1 2956
box -32 -32 32 32
use via_M1_M2_1_l  NoName_214 ~/A2G/MAGIC/magic_layout/skywater130_microtemplates_dense
timestamp 1647525606
transform 1 0 3438 0 1 2444
box -32 -32 32 32
use via_M1_M2_1_m  NoName_215 ~/A2G/MAGIC/magic_layout/skywater130_microtemplates_dense
timestamp 1647525606
transform 1 0 3438 0 1 3084
box -32 -32 32 32
use via_M1_M2_1_n  NoName_216 ~/A2G/MAGIC/magic_layout/skywater130_microtemplates_dense
timestamp 1647525606
transform 1 0 3438 0 1 2316
box -32 -32 32 32
use via_M1_M2_1_o  NoName_217 ~/A2G/MAGIC/magic_layout/skywater130_microtemplates_dense
timestamp 1647525606
transform 1 0 6762 0 1 900
box -32 -32 32 32
use via_M1_M2_1_p  NoName_218 ~/A2G/MAGIC/magic_layout/skywater130_microtemplates_dense
timestamp 1647525606
transform 1 0 6762 0 1 1028
box -32 -32 32 32
use via_M1_M2_1_q  NoName_219 ~/A2G/MAGIC/magic_layout/skywater130_microtemplates_dense
timestamp 1647525606
transform 1 0 6762 0 1 772
box -32 -32 32 32
use via_M1_M2_1_r  NoName_220 ~/A2G/MAGIC/magic_layout/skywater130_microtemplates_dense
timestamp 1647525606
transform 1 0 6762 0 1 1156
box -32 -32 32 32
use via_M1_M2_1_s  NoName_221 ~/A2G/MAGIC/magic_layout/skywater130_microtemplates_dense
timestamp 1647525606
transform 1 0 6762 0 1 644
box -32 -32 32 32
use via_M1_M2_1_t  NoName_222 ~/A2G/MAGIC/magic_layout/skywater130_microtemplates_dense
timestamp 1647525606
transform 1 0 6762 0 1 1284
box -32 -32 32 32
use via_M1_M2_1_u  NoName_223 ~/A2G/MAGIC/magic_layout/skywater130_microtemplates_dense
timestamp 1647525606
transform 1 0 6762 0 1 516
box -32 -32 32 32
use via_M1_M2_1_v  NoName_224 ~/A2G/MAGIC/magic_layout/skywater130_microtemplates_dense
timestamp 1647525606
transform 1 0 9038 0 1 900
box -32 -32 32 32
use via_M1_M2_1_w  NoName_225 ~/A2G/MAGIC/magic_layout/skywater130_microtemplates_dense
timestamp 1647525606
transform 1 0 9038 0 1 1028
box -32 -32 32 32
use via_M1_M2_1_x  NoName_226 ~/A2G/MAGIC/magic_layout/skywater130_microtemplates_dense
timestamp 1647525606
transform 1 0 9038 0 1 772
box -32 -32 32 32
use via_M1_M2_1_y  NoName_227 ~/A2G/MAGIC/magic_layout/skywater130_microtemplates_dense
timestamp 1647525606
transform 1 0 9038 0 1 1156
box -32 -32 32 32
use via_M1_M2_1_z  NoName_228 ~/A2G/MAGIC/magic_layout/skywater130_microtemplates_dense
timestamp 1647525606
transform 1 0 9038 0 1 644
box -32 -32 32 32
use via_M1_M2_1_{  NoName_229 ~/A2G/MAGIC/magic_layout/skywater130_microtemplates_dense
timestamp 1647525606
transform 1 0 9038 0 1 1284
box -32 -32 32 32
use via_M1_M2_1_|  NoName_230 ~/A2G/MAGIC/magic_layout/skywater130_microtemplates_dense
timestamp 1647525606
transform 1 0 9038 0 1 516
box -32 -32 32 32
use via_M1_M2_1_}  NoName_231 ~/A2G/MAGIC/magic_layout/skywater130_microtemplates_dense
timestamp 1647525606
transform 1 0 6762 0 1 2700
box -32 -32 32 32
use via_M1_M2_1_~  NoName_232 ~/A2G/MAGIC/magic_layout/skywater130_microtemplates_dense
timestamp 1647525606
transform 1 0 6762 0 1 2828
box -32 -32 32 32
use via_M1_M2_1_  NoName_233 ~/A2G/MAGIC/magic_layout/skywater130_microtemplates_dense
timestamp 1647525606
transform 1 0 6762 0 1 2572
box -32 -32 32 32
use via_M1_M2_1_�  NoName_234 ~/A2G/MAGIC/magic_layout/skywater130_microtemplates_dense
timestamp 1647525606
transform 1 0 6762 0 1 2956
box -32 -32 32 32
use via_M1_M2_1_�  NoName_235 ~/A2G/MAGIC/magic_layout/skywater130_microtemplates_dense
timestamp 1647525606
transform 1 0 6762 0 1 2444
box -32 -32 32 32
use via_M1_M2_1_�  NoName_236 ~/A2G/MAGIC/magic_layout/skywater130_microtemplates_dense
timestamp 1647525606
transform 1 0 6762 0 1 3084
box -32 -32 32 32
use via_M1_M2_1_�  NoName_237 ~/A2G/MAGIC/magic_layout/skywater130_microtemplates_dense
timestamp 1647525606
transform 1 0 6762 0 1 2316
box -32 -32 32 32
use via_M1_M2_1_�  NoName_238 ~/A2G/MAGIC/magic_layout/skywater130_microtemplates_dense
timestamp 1647525606
transform 1 0 9038 0 1 2700
box -32 -32 32 32
use via_M1_M2_1_�  NoName_239 ~/A2G/MAGIC/magic_layout/skywater130_microtemplates_dense
timestamp 1647525606
transform 1 0 9038 0 1 2828
box -32 -32 32 32
use via_M1_M2_1_�  NoName_240 ~/A2G/MAGIC/magic_layout/skywater130_microtemplates_dense
timestamp 1647525606
transform 1 0 9038 0 1 2572
box -32 -32 32 32
use via_M1_M2_1_�  NoName_241 ~/A2G/MAGIC/magic_layout/skywater130_microtemplates_dense
timestamp 1647525606
transform 1 0 9038 0 1 2956
box -32 -32 32 32
use via_M1_M2_1_�  NoName_242 ~/A2G/MAGIC/magic_layout/skywater130_microtemplates_dense
timestamp 1647525606
transform 1 0 9038 0 1 2444
box -32 -32 32 32
use via_M1_M2_1_�  NoName_243 ~/A2G/MAGIC/magic_layout/skywater130_microtemplates_dense
timestamp 1647525606
transform 1 0 9038 0 1 3084
box -32 -32 32 32
use via_M1_M2_1_�  NoName_244 ~/A2G/MAGIC/magic_layout/skywater130_microtemplates_dense
timestamp 1647525606
transform 1 0 9038 0 1 2316
box -32 -32 32 32
use via_M1_M2_1_�  NoName_245 ~/A2G/MAGIC/magic_layout/skywater130_microtemplates_dense
timestamp 1647525606
transform 1 0 1162 0 1 900
box -32 -32 32 32
use via_M1_M2_1_�  NoName_246 ~/A2G/MAGIC/magic_layout/skywater130_microtemplates_dense
timestamp 1647525606
transform 1 0 1162 0 1 1028
box -32 -32 32 32
use via_M1_M2_1_�  NoName_247 ~/A2G/MAGIC/magic_layout/skywater130_microtemplates_dense
timestamp 1647525606
transform 1 0 1162 0 1 772
box -32 -32 32 32
use via_M1_M2_1_�  NoName_248 ~/A2G/MAGIC/magic_layout/skywater130_microtemplates_dense
timestamp 1647525606
transform 1 0 1162 0 1 1156
box -32 -32 32 32
use via_M1_M2_1_�  NoName_249 ~/A2G/MAGIC/magic_layout/skywater130_microtemplates_dense
timestamp 1647525606
transform 1 0 1162 0 1 644
box -32 -32 32 32
use via_M1_M2_1_�  NoName_250 ~/A2G/MAGIC/magic_layout/skywater130_microtemplates_dense
timestamp 1647525606
transform 1 0 1162 0 1 1284
box -32 -32 32 32
use via_M1_M2_1_�  NoName_251 ~/A2G/MAGIC/magic_layout/skywater130_microtemplates_dense
timestamp 1647525606
transform 1 0 1162 0 1 516
box -32 -32 32 32
use via_M1_M2_1_�  NoName_252 ~/A2G/MAGIC/magic_layout/skywater130_microtemplates_dense
timestamp 1647525606
transform 1 0 3438 0 1 900
box -32 -32 32 32
use via_M1_M2_1_�  NoName_253 ~/A2G/MAGIC/magic_layout/skywater130_microtemplates_dense
timestamp 1647525606
transform 1 0 3438 0 1 1028
box -32 -32 32 32
use via_M1_M2_1_�  NoName_254 ~/A2G/MAGIC/magic_layout/skywater130_microtemplates_dense
timestamp 1647525606
transform 1 0 3438 0 1 772
box -32 -32 32 32
use via_M1_M2_1_�  NoName_255 ~/A2G/MAGIC/magic_layout/skywater130_microtemplates_dense
timestamp 1647525606
transform 1 0 3438 0 1 1156
box -32 -32 32 32
use via_M1_M2_1_�  NoName_256 ~/A2G/MAGIC/magic_layout/skywater130_microtemplates_dense
timestamp 1647525606
transform 1 0 3438 0 1 644
box -32 -32 32 32
use via_M1_M2_1_�  NoName_257 ~/A2G/MAGIC/magic_layout/skywater130_microtemplates_dense
timestamp 1647525606
transform 1 0 3438 0 1 1284
box -32 -32 32 32
use via_M1_M2_1_�  NoName_258 ~/A2G/MAGIC/magic_layout/skywater130_microtemplates_dense
timestamp 1647525606
transform 1 0 3438 0 1 516
box -32 -32 32 32
use via_M1_M2_1_�  NoName_259 ~/A2G/MAGIC/magic_layout/skywater130_microtemplates_dense
timestamp 1647525606
transform 1 0 3960 0 1 2700
box -32 -32 32 32
use via_M1_M2_1_�  NoName_260 ~/A2G/MAGIC/magic_layout/skywater130_microtemplates_dense
timestamp 1647525606
transform 1 0 3960 0 1 2828
box -32 -32 32 32
use via_M1_M2_1_�  NoName_261 ~/A2G/MAGIC/magic_layout/skywater130_microtemplates_dense
timestamp 1647525606
transform 1 0 3960 0 1 2572
box -32 -32 32 32
use via_M1_M2_1_�  NoName_262 ~/A2G/MAGIC/magic_layout/skywater130_microtemplates_dense
timestamp 1647525606
transform 1 0 3960 0 1 2956
box -32 -32 32 32
use via_M1_M2_1_�  NoName_263 ~/A2G/MAGIC/magic_layout/skywater130_microtemplates_dense
timestamp 1647525606
transform 1 0 3960 0 1 2444
box -32 -32 32 32
use via_M1_M2_1_�  NoName_264 ~/A2G/MAGIC/magic_layout/skywater130_microtemplates_dense
timestamp 1647525606
transform 1 0 3960 0 1 3084
box -32 -32 32 32
use via_M1_M2_1_�  NoName_265 ~/A2G/MAGIC/magic_layout/skywater130_microtemplates_dense
timestamp 1647525606
transform 1 0 3960 0 1 2316
box -32 -32 32 32
use via_M1_M2_1_�  NoName_266 ~/A2G/MAGIC/magic_layout/skywater130_microtemplates_dense
timestamp 1647525606
transform 1 0 6238 0 1 2700
box -32 -32 32 32
use via_M1_M2_1_�  NoName_267 ~/A2G/MAGIC/magic_layout/skywater130_microtemplates_dense
timestamp 1647525606
transform 1 0 6238 0 1 2828
box -32 -32 32 32
use via_M1_M2_1_�  NoName_268 ~/A2G/MAGIC/magic_layout/skywater130_microtemplates_dense
timestamp 1647525606
transform 1 0 6238 0 1 2572
box -32 -32 32 32
use via_M1_M2_1_�  NoName_269 ~/A2G/MAGIC/magic_layout/skywater130_microtemplates_dense
timestamp 1647525606
transform 1 0 6238 0 1 2956
box -32 -32 32 32
use via_M1_M2_1_�  NoName_270 ~/A2G/MAGIC/magic_layout/skywater130_microtemplates_dense
timestamp 1647525606
transform 1 0 6238 0 1 2444
box -32 -32 32 32
use via_M1_M2_1_�  NoName_271 ~/A2G/MAGIC/magic_layout/skywater130_microtemplates_dense
timestamp 1647525606
transform 1 0 6238 0 1 3084
box -32 -32 32 32
use via_M1_M2_1_�  NoName_272 ~/A2G/MAGIC/magic_layout/skywater130_microtemplates_dense
timestamp 1647525606
transform 1 0 6238 0 1 2316
box -32 -32 32 32
use via_M1_M2_1_�  NoName_273 ~/A2G/MAGIC/magic_layout/skywater130_microtemplates_dense
timestamp 1647525606
transform 1 0 3960 0 1 900
box -32 -32 32 32
use via_M1_M2_1_�  NoName_274 ~/A2G/MAGIC/magic_layout/skywater130_microtemplates_dense
timestamp 1647525606
transform 1 0 3960 0 1 1028
box -32 -32 32 32
use via_M1_M2_1_�  NoName_275 ~/A2G/MAGIC/magic_layout/skywater130_microtemplates_dense
timestamp 1647525606
transform 1 0 3960 0 1 772
box -32 -32 32 32
use via_M1_M2_1_�  NoName_276 ~/A2G/MAGIC/magic_layout/skywater130_microtemplates_dense
timestamp 1647525606
transform 1 0 3960 0 1 1156
box -32 -32 32 32
use via_M1_M2_1_�  NoName_277 ~/A2G/MAGIC/magic_layout/skywater130_microtemplates_dense
timestamp 1647525606
transform 1 0 3960 0 1 644
box -32 -32 32 32
use via_M1_M2_1_�  NoName_278 ~/A2G/MAGIC/magic_layout/skywater130_microtemplates_dense
timestamp 1647525606
transform 1 0 3960 0 1 1284
box -32 -32 32 32
use via_M1_M2_1_�  NoName_279 ~/A2G/MAGIC/magic_layout/skywater130_microtemplates_dense
timestamp 1647525606
transform 1 0 3960 0 1 516
box -32 -32 32 32
use via_M1_M2_1_�  NoName_280 ~/A2G/MAGIC/magic_layout/skywater130_microtemplates_dense
timestamp 1647525606
transform 1 0 6238 0 1 900
box -32 -32 32 32
use via_M1_M2_1_�  NoName_281 ~/A2G/MAGIC/magic_layout/skywater130_microtemplates_dense
timestamp 1647525606
transform 1 0 6238 0 1 1028
box -32 -32 32 32
use via_M1_M2_1_�  NoName_282 ~/A2G/MAGIC/magic_layout/skywater130_microtemplates_dense
timestamp 1647525606
transform 1 0 6238 0 1 772
box -32 -32 32 32
use via_M1_M2_1_�  NoName_283 ~/A2G/MAGIC/magic_layout/skywater130_microtemplates_dense
timestamp 1647525606
transform 1 0 6238 0 1 1156
box -32 -32 32 32
use via_M1_M2_1_�  NoName_284 ~/A2G/MAGIC/magic_layout/skywater130_microtemplates_dense
timestamp 1647525606
transform 1 0 6238 0 1 644
box -32 -32 32 32
use via_M1_M2_1_�  NoName_285 ~/A2G/MAGIC/magic_layout/skywater130_microtemplates_dense
timestamp 1647525606
transform 1 0 6238 0 1 1284
box -32 -32 32 32
use via_M1_M2_1_�  NoName_286 ~/A2G/MAGIC/magic_layout/skywater130_microtemplates_dense
timestamp 1647525606
transform 1 0 6238 0 1 516
box -32 -32 32 32
use via_M2_M3_0  NoName_287 ~/A2G/MAGIC/magic_layout/skywater130_microtemplates_dense
timestamp 1647525786
transform 1 0 2300 0 1 2700
box -38 -38 38 38
use via_M2_M3_0  NoName_288
timestamp 1647525786
transform 1 0 2300 0 1 900
box -38 -38 38 38
use via_M2_M3_0  NoName_291
timestamp 1647525786
transform 1 0 7900 0 1 900
box -38 -38 38 38
use via_M2_M3_0  NoName_292
timestamp 1647525786
transform 1 0 7900 0 1 2700
box -38 -38 38 38
use via_M2_M3_0  NoName_295
timestamp 1647525786
transform 1 0 3100 0 1 500
box -38 -38 38 38
use via_M2_M3_0  NoName_296
timestamp 1647525786
transform 1 0 4100 0 1 900
box -38 -38 38 38
use via_M2_M3_0  NoName_299
timestamp 1647525786
transform 1 0 7100 0 1 500
box -38 -38 38 38
use via_M2_M3_0  NoName_300
timestamp 1647525786
transform 1 0 6100 0 1 900
box -38 -38 38 38
use via_M2_M3_0  NoName_303
timestamp 1647525786
transform 1 0 1300 0 1 900
box -38 -38 38 38
use via_M2_M3_0  NoName_305
timestamp 1647525786
transform 1 0 500 0 1 900
box -38 -38 38 38
use via_M2_M3_0  NoName_306
timestamp 1647525786
transform 1 0 8900 0 1 900
box -38 -38 38 38
use via_M2_M3_0  NoName_308
timestamp 1647525786
transform 1 0 9700 0 1 900
box -38 -38 38 38
use via_M2_M3_0  NoName_309
timestamp 1647525786
transform 1 0 3300 0 1 900
box -38 -38 38 38
use via_M2_M3_0  NoName_310
timestamp 1647525786
transform 1 0 7100 0 1 1300
box -38 -38 38 38
use via_M2_M3_0  NoName_313
timestamp 1647525786
transform 1 0 6900 0 1 900
box -38 -38 38 38
use via_M2_M3_0  NoName_314
timestamp 1647525786
transform 1 0 3100 0 1 1300
box -38 -38 38 38
use via_M3_M4_0  NoName_316 ~/A2G/MAGIC/magic_layout/skywater130_microtemplates_dense
timestamp 1647526059
transform 1 0 6700 0 1 900
box -38 -38 38 38
use via_M3_M4_0  NoName_317
timestamp 1647526059
transform 1 0 3100 0 1 1100
box -38 -38 38 38
use via_M2_M3_0  NoName_319
timestamp 1647525786
transform 1 0 3100 0 1 2300
box -38 -38 38 38
use via_M2_M3_0  NoName_320
timestamp 1647525786
transform 1 0 4100 0 1 2700
box -38 -38 38 38
use via_M2_M3_0  NoName_323
timestamp 1647525786
transform 1 0 7100 0 1 2300
box -38 -38 38 38
use via_M2_M3_0  NoName_324
timestamp 1647525786
transform 1 0 6100 0 1 2700
box -38 -38 38 38
use via_M1_M2_1_�  NoName_327 ~/A2G/MAGIC/magic_layout/skywater130_microtemplates_dense
timestamp 1647525606
transform 1 0 500 0 1 2750
box -32 -32 32 32
use via_M1_M2_1_�  NoName_328 ~/A2G/MAGIC/magic_layout/skywater130_microtemplates_dense
timestamp 1647525606
transform 1 0 9700 0 1 2750
box -32 -32 32 32
use XM1  XM1 ~/A2G/MAGIC/magic_layout/pcell
timestamp 1679988681
transform 1 0 2300 0 1 2700
box -1191 -529 1191 529
use XM2  XM2 ~/A2G/MAGIC/magic_layout/pcell
timestamp 1679988681
transform -1 0 7900 0 -1 900
box -1191 -529 1191 529
use XM3  XM3 ~/A2G/MAGIC/magic_layout/pcell
timestamp 1679988682
transform 1 0 7900 0 1 2700
box -1191 -529 1191 529
use XM4  XM4 ~/A2G/MAGIC/magic_layout/pcell
timestamp 1679988682
transform -1 0 2300 0 -1 900
box -1191 -529 1191 529
use XM5  XM5 ~/A2G/MAGIC/magic_layout/pcell
timestamp 1679988683
transform 1 0 5100 0 1 2700
box -1191 -529 1191 529
use XM6  XM6 ~/A2G/MAGIC/magic_layout/pcell
timestamp 1679988683
transform -1 0 5100 0 -1 900
box -1191 -529 1191 529
use XR1  XR1 ~/A2G/MAGIC/magic_layout/pcell
timestamp 1679988684
transform -1 0 500 0 -1 1700
box -258 -1061 258 1061
use XR2  XR2 ~/A2G/MAGIC/magic_layout/pcell
timestamp 1679988684
transform -1 0 9700 0 -1 1700
box -258 -1061 258 1061
<< labels >>
flabel metal3 5100 1300 5100 1300 0 FreeSans 1600 0 0 0 oa
flabel metal4 4900 1100 4900 1100 0 FreeSans 1600 0 0 0 ob
flabel metal2 2300 3100 2300 3100 0 FreeSans 1600 0 0 0 ia
flabel metal2 7900 3100 7900 3100 0 FreeSans 1600 0 0 0 ib
flabel metal2 5100 3100 5100 3100 0 FreeSans 1600 0 0 0 icmlbias
flabel metal2 5100 500 5100 500 0 FreeSans 1600 0 0 0 ihysbias
flabel metal2 500 2500 500 2500 0 FreeSans 1600 0 0 0 vdd
flabel metal2 9700 2500 9700 2500 0 FreeSans 1600 0 0 0 vdd
flabel metal2 5100 2300 5100 2300 0 FreeSans 1600 0 0 0 vss
flabel metal2 5100 1290 5100 1290 0 FreeSans 1600 0 0 0 vss
<< end >>
