* NGSPICE file created from diff2sin.ext - technology: sky130A

.subckt XM1_origin G D S a_n1155_n493#
X0 S G D a_n1155_n493# sky130_fd_pr__nfet_01v8_lvt ad=8.12e+12p pd=6.064e+07u as=9.135e+12p ps=6.822e+07u w=3.5e+06u l=350000u
X1 S G D a_n1155_n493# sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=3.5e+06u l=350000u
X2 S G D a_n1155_n493# sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=3.5e+06u l=350000u
X3 D G S a_n1155_n493# sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=3.5e+06u l=350000u
X4 D G S a_n1155_n493# sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=3.5e+06u l=350000u
X5 S G D a_n1155_n493# sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=3.5e+06u l=350000u
X6 D G S a_n1155_n493# sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=3.5e+06u l=350000u
X7 S G D a_n1155_n493# sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=3.5e+06u l=350000u
X8 D G S a_n1155_n493# sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=3.5e+06u l=350000u
X9 S G D a_n1155_n493# sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=3.5e+06u l=350000u
X10 S G D a_n1155_n493# sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=3.5e+06u l=350000u
X11 S G D a_n1155_n493# sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=3.5e+06u l=350000u
X12 D G S a_n1155_n493# sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=3.5e+06u l=350000u
X13 D G S a_n1155_n493# sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=3.5e+06u l=350000u
X14 D G S a_n1155_n493# sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=3.5e+06u l=350000u
X15 D G S a_n1155_n493# sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=3.5e+06u l=350000u
C0 S D 10.12fF
C1 D a_n1155_n493# 0.86fF
C2 S a_n1155_n493# 0.37fF
C3 G a_n1155_n493# 3.39fF
.ends

.subckt XM1 XM1/S XM1/G XM1/D VSUBS
XXM1 XM1/G XM1/D XM1/S VSUBS XM1_origin
C0 XM1/G XM1/S 0.57fF
C1 XM1/G XM1/D 1.19fF
C2 XM1/D XM1/S 1.24fF
C3 XM1/D VSUBS 0.91fF
C4 XM1/G VSUBS 4.45fF
C5 XM1/S VSUBS 0.93fF
.ends

.subckt XM2_origin G D S w_n2727_n534# VSUBS
X0 S G D w_n2727_n534# sky130_fd_pr__pfet_01v8_lvt ad=2.03e+13p pd=1.516e+08u as=2.1315e+13p ps=1.5918e+08u w=3.5e+06u l=350000u
X1 D G S w_n2727_n534# sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=3.5e+06u l=350000u
X2 D G S w_n2727_n534# sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=3.5e+06u l=350000u
X3 D G S w_n2727_n534# sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=3.5e+06u l=350000u
X4 S G D w_n2727_n534# sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=3.5e+06u l=350000u
X5 S G D w_n2727_n534# sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=3.5e+06u l=350000u
X6 S G D w_n2727_n534# sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=3.5e+06u l=350000u
X7 S G D w_n2727_n534# sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=3.5e+06u l=350000u
X8 S G D w_n2727_n534# sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=3.5e+06u l=350000u
X9 S G D w_n2727_n534# sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=3.5e+06u l=350000u
X10 D G S w_n2727_n534# sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=3.5e+06u l=350000u
X11 D G S w_n2727_n534# sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=3.5e+06u l=350000u
X12 D G S w_n2727_n534# sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=3.5e+06u l=350000u
X13 D G S w_n2727_n534# sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=3.5e+06u l=350000u
X14 S G D w_n2727_n534# sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=3.5e+06u l=350000u
X15 S G D w_n2727_n534# sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=3.5e+06u l=350000u
X16 S G D w_n2727_n534# sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=3.5e+06u l=350000u
X17 S G D w_n2727_n534# sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=3.5e+06u l=350000u
X18 D G S w_n2727_n534# sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=3.5e+06u l=350000u
X19 D G S w_n2727_n534# sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=3.5e+06u l=350000u
X20 D G S w_n2727_n534# sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=3.5e+06u l=350000u
X21 D G S w_n2727_n534# sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=3.5e+06u l=350000u
X22 D G S w_n2727_n534# sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=3.5e+06u l=350000u
X23 D G S w_n2727_n534# sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=3.5e+06u l=350000u
X24 S G D w_n2727_n534# sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=3.5e+06u l=350000u
X25 S G D w_n2727_n534# sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=3.5e+06u l=350000u
X26 S G D w_n2727_n534# sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=3.5e+06u l=350000u
X27 S G D w_n2727_n534# sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=3.5e+06u l=350000u
X28 S G D w_n2727_n534# sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=3.5e+06u l=350000u
X29 S G D w_n2727_n534# sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=3.5e+06u l=350000u
X30 D G S w_n2727_n534# sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=3.5e+06u l=350000u
X31 D G S w_n2727_n534# sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=3.5e+06u l=350000u
X32 D G S w_n2727_n534# sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=3.5e+06u l=350000u
X33 D G S w_n2727_n534# sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=3.5e+06u l=350000u
X34 D G S w_n2727_n534# sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=3.5e+06u l=350000u
X35 D G S w_n2727_n534# sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=3.5e+06u l=350000u
X36 D G S w_n2727_n534# sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=3.5e+06u l=350000u
X37 S G D w_n2727_n534# sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=3.5e+06u l=350000u
X38 S G D w_n2727_n534# sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=3.5e+06u l=350000u
X39 S G D w_n2727_n534# sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=3.5e+06u l=350000u
C0 D w_n2727_n534# 1.39fF
C1 D S 25.31fF
C2 w_n2727_n534# G 7.77fF
C3 w_n2727_n534# S 0.90fF
C4 G VSUBS 0.91fF
C5 w_n2727_n534# VSUBS 17.47fF
.ends

.subckt XM2 XM2/w_n2727_n534# XM2/S XM2/G XM2/D VSUBS
XXM2 XM2/G XM2/D XM2/S XM2/w_n2727_n534# VSUBS XM2_origin
C0 XM2/S XM2/D 3.31fF
C1 XM2/S XM2/w_n2727_n534# 1.40fF
C2 XM2/D XM2/w_n2727_n534# 0.06fF
C3 XM2/G XM2/S 1.52fF
C4 XM2/G XM2/D 3.01fF
C5 XM2/G XM2/w_n2727_n534# 2.59fF
C6 XM2/w_n2727_n534# VSUBS 17.47fF
C7 XM2/G VSUBS 0.91fF
.ends

.subckt XM3_origin G D S a_n1155_n493#
X0 S G D a_n1155_n493# sky130_fd_pr__nfet_01v8_lvt ad=8.12e+12p pd=6.064e+07u as=9.135e+12p ps=6.822e+07u w=3.5e+06u l=350000u
X1 S G D a_n1155_n493# sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=3.5e+06u l=350000u
X2 S G D a_n1155_n493# sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=3.5e+06u l=350000u
X3 D G S a_n1155_n493# sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=3.5e+06u l=350000u
X4 D G S a_n1155_n493# sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=3.5e+06u l=350000u
X5 S G D a_n1155_n493# sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=3.5e+06u l=350000u
X6 D G S a_n1155_n493# sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=3.5e+06u l=350000u
X7 S G D a_n1155_n493# sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=3.5e+06u l=350000u
X8 D G S a_n1155_n493# sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=3.5e+06u l=350000u
X9 S G D a_n1155_n493# sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=3.5e+06u l=350000u
X10 S G D a_n1155_n493# sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=3.5e+06u l=350000u
X11 S G D a_n1155_n493# sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=3.5e+06u l=350000u
X12 D G S a_n1155_n493# sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=3.5e+06u l=350000u
X13 D G S a_n1155_n493# sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=3.5e+06u l=350000u
X14 D G S a_n1155_n493# sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=3.5e+06u l=350000u
X15 D G S a_n1155_n493# sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=3.5e+06u l=350000u
C0 D S 10.12fF
C1 D a_n1155_n493# 0.86fF
C2 S a_n1155_n493# 0.37fF
C3 G a_n1155_n493# 3.39fF
.ends

.subckt XM3 XM3/D XM3/S XM3/G VSUBS
XXM3 XM3/G XM3/D XM3/S VSUBS XM3_origin
C0 XM3/S XM3/D 1.24fF
C1 XM3/G XM3/D 1.19fF
C2 XM3/G XM3/S 0.57fF
C3 XM3/D VSUBS 0.91fF
C4 XM3/S VSUBS 0.93fF
C5 XM3/G VSUBS 4.45fF
.ends

.subckt XM4_origin G D S w_n2727_n534# VSUBS
X0 S G D w_n2727_n534# sky130_fd_pr__pfet_01v8_lvt ad=2.03e+13p pd=1.516e+08u as=2.1315e+13p ps=1.5918e+08u w=3.5e+06u l=350000u
X1 D G S w_n2727_n534# sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=3.5e+06u l=350000u
X2 D G S w_n2727_n534# sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=3.5e+06u l=350000u
X3 D G S w_n2727_n534# sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=3.5e+06u l=350000u
X4 S G D w_n2727_n534# sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=3.5e+06u l=350000u
X5 S G D w_n2727_n534# sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=3.5e+06u l=350000u
X6 S G D w_n2727_n534# sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=3.5e+06u l=350000u
X7 S G D w_n2727_n534# sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=3.5e+06u l=350000u
X8 S G D w_n2727_n534# sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=3.5e+06u l=350000u
X9 S G D w_n2727_n534# sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=3.5e+06u l=350000u
X10 D G S w_n2727_n534# sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=3.5e+06u l=350000u
X11 D G S w_n2727_n534# sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=3.5e+06u l=350000u
X12 D G S w_n2727_n534# sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=3.5e+06u l=350000u
X13 D G S w_n2727_n534# sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=3.5e+06u l=350000u
X14 S G D w_n2727_n534# sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=3.5e+06u l=350000u
X15 S G D w_n2727_n534# sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=3.5e+06u l=350000u
X16 S G D w_n2727_n534# sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=3.5e+06u l=350000u
X17 S G D w_n2727_n534# sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=3.5e+06u l=350000u
X18 D G S w_n2727_n534# sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=3.5e+06u l=350000u
X19 D G S w_n2727_n534# sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=3.5e+06u l=350000u
X20 D G S w_n2727_n534# sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=3.5e+06u l=350000u
X21 D G S w_n2727_n534# sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=3.5e+06u l=350000u
X22 D G S w_n2727_n534# sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=3.5e+06u l=350000u
X23 D G S w_n2727_n534# sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=3.5e+06u l=350000u
X24 S G D w_n2727_n534# sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=3.5e+06u l=350000u
X25 S G D w_n2727_n534# sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=3.5e+06u l=350000u
X26 S G D w_n2727_n534# sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=3.5e+06u l=350000u
X27 S G D w_n2727_n534# sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=3.5e+06u l=350000u
X28 S G D w_n2727_n534# sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=3.5e+06u l=350000u
X29 S G D w_n2727_n534# sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=3.5e+06u l=350000u
X30 D G S w_n2727_n534# sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=3.5e+06u l=350000u
X31 D G S w_n2727_n534# sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=3.5e+06u l=350000u
X32 D G S w_n2727_n534# sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=3.5e+06u l=350000u
X33 D G S w_n2727_n534# sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=3.5e+06u l=350000u
X34 D G S w_n2727_n534# sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=3.5e+06u l=350000u
X35 D G S w_n2727_n534# sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=3.5e+06u l=350000u
X36 D G S w_n2727_n534# sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=3.5e+06u l=350000u
X37 S G D w_n2727_n534# sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=3.5e+06u l=350000u
X38 S G D w_n2727_n534# sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=3.5e+06u l=350000u
X39 S G D w_n2727_n534# sky130_fd_pr__pfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=3.5e+06u l=350000u
C0 S D 25.31fF
C1 w_n2727_n534# S 0.90fF
C2 w_n2727_n534# D 1.39fF
C3 w_n2727_n534# G 7.77fF
C4 G VSUBS 0.91fF
C5 w_n2727_n534# VSUBS 17.47fF
.ends

.subckt XM4 XM4/S XM4/G XM4/D XM4/w_n2727_n534# VSUBS
XXM4 XM4/G XM4/D XM4/S XM4/w_n2727_n534# VSUBS XM4_origin
C0 XM4/D XM4/S 3.31fF
C1 XM4/G XM4/w_n2727_n534# 2.59fF
C2 XM4/S XM4/w_n2727_n534# 1.40fF
C3 XM4/D XM4/w_n2727_n534# 0.06fF
C4 XM4/G XM4/S 1.52fF
C5 XM4/G XM4/D 3.01fF
C6 XM4/G VSUBS 0.91fF
C7 XM4/w_n2727_n534# VSUBS 17.47fF
.ends

.subckt XM5_origin G D S a_n2179_n493#
X0 S G D a_n2179_n493# sky130_fd_pr__nfet_01v8_lvt ad=1.624e+13p pd=1.2128e+08u as=1.7255e+13p ps=1.2886e+08u w=3.5e+06u l=350000u
X1 S G D a_n2179_n493# sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=3.5e+06u l=350000u
X2 S G D a_n2179_n493# sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=3.5e+06u l=350000u
X3 S G D a_n2179_n493# sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=3.5e+06u l=350000u
X4 S G D a_n2179_n493# sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=3.5e+06u l=350000u
X5 D G S a_n2179_n493# sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=3.5e+06u l=350000u
X6 D G S a_n2179_n493# sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=3.5e+06u l=350000u
X7 D G S a_n2179_n493# sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=3.5e+06u l=350000u
X8 D G S a_n2179_n493# sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=3.5e+06u l=350000u
X9 D G S a_n2179_n493# sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=3.5e+06u l=350000u
X10 S G D a_n2179_n493# sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=3.5e+06u l=350000u
X11 D G S a_n2179_n493# sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=3.5e+06u l=350000u
X12 S G D a_n2179_n493# sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=3.5e+06u l=350000u
X13 S G D a_n2179_n493# sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=3.5e+06u l=350000u
X14 D G S a_n2179_n493# sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=3.5e+06u l=350000u
X15 D G S a_n2179_n493# sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=3.5e+06u l=350000u
X16 D G S a_n2179_n493# sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=3.5e+06u l=350000u
X17 S G D a_n2179_n493# sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=3.5e+06u l=350000u
X18 S G D a_n2179_n493# sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=3.5e+06u l=350000u
X19 S G D a_n2179_n493# sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=3.5e+06u l=350000u
X20 S G D a_n2179_n493# sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=3.5e+06u l=350000u
X21 S G D a_n2179_n493# sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=3.5e+06u l=350000u
X22 D G S a_n2179_n493# sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=3.5e+06u l=350000u
X23 D G S a_n2179_n493# sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=3.5e+06u l=350000u
X24 S G D a_n2179_n493# sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=3.5e+06u l=350000u
X25 S G D a_n2179_n493# sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=3.5e+06u l=350000u
X26 S G D a_n2179_n493# sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=3.5e+06u l=350000u
X27 D G S a_n2179_n493# sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=3.5e+06u l=350000u
X28 D G S a_n2179_n493# sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=3.5e+06u l=350000u
X29 D G S a_n2179_n493# sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=3.5e+06u l=350000u
X30 D G S a_n2179_n493# sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=3.5e+06u l=350000u
X31 D G S a_n2179_n493# sky130_fd_pr__nfet_01v8_lvt ad=0p pd=0u as=0p ps=0u w=3.5e+06u l=350000u
C0 S D 20.25fF
C1 D a_n2179_n493# 1.22fF
C2 S a_n2179_n493# 0.73fF
C3 G a_n2179_n493# 6.75fF
.ends

.subckt XM5 XM5/G XM5/D XM5/S VSUBS
XXM5 XM5/G XM5/D XM5/S VSUBS XM5_origin
C0 XM5/D XM5/S 2.57fF
C1 XM5/G XM5/S 1.17fF
C2 XM5/D XM5/G 2.40fF
C3 XM5/D VSUBS 1.28fF
C4 XM5/S VSUBS 1.89fF
C5 XM5/G VSUBS 8.88fF
.ends

.subckt diff2sin out ia ib icmbias vdd vss
XXM1 XM5/XM5/D ia XM4/XM4/G vss XM1
XXM2 vdd vdd XM4/XM4/G XM4/XM4/G vss XM2
XXM3 out XM5/XM5/D ib vss XM3
XXM4 vdd XM4/XM4/G out vdd vss XM4
XXM5 icmbias XM5/XM5/D vss vss XM5
C0 vdd XM4/XM4/G 3.12fF
C1 out ib 0.34fF
C2 XM5/XM5/D out 0.53fF
C3 XM5/XM5/D ib 0.25fF
C4 vdd out 1.48fF
C5 ia XM5/XM5/D 0.25fF
C6 XM5/XM5/D icmbias 0.15fF
C7 vdd ib 0.19fF
C8 vdd ia 0.19fF
C9 vdd icmbias 0.40fF
C10 vdd XM5/XM5/D 0.43fF
C11 XM4/XM4/G out 0.30fF
C12 ia XM4/XM4/G 0.34fF
C13 XM5/XM5/D XM4/XM4/G 0.53fF
C14 XM5/XM5/D vss 6.48fF
C15 icmbias vss 9.90fF
C16 out vss 2.52fF
C17 ib vss 5.00fF
C18 vdd vss 135.37fF
C19 XM4/XM4/G vss 7.27fF
C20 ia vss 5.00fF
.ends

